  --Example instantiation for system 'nios2_fpu'
  nios2_fpu_inst : nios2_fpu
    port map(
      AUD_L_from_the_spu => AUD_L_from_the_spu,
      AUD_R_from_the_spu => AUD_R_from_the_spu,
      DAC_BCLK_from_the_spu => DAC_BCLK_from_the_spu,
      DAC_DATA_from_the_spu => DAC_DATA_from_the_spu,
      DAC_LRCK_from_the_spu => DAC_LRCK_from_the_spu,
      MMC_SCK_from_the_mmcdma => MMC_SCK_from_the_mmcdma,
      MMC_SDO_from_the_mmcdma => MMC_SDO_from_the_mmcdma,
      MMC_nCS_from_the_mmcdma => MMC_nCS_from_the_mmcdma,
      PS2_CLK_to_and_from_the_ps2_keyboard => PS2_CLK_to_and_from_the_ps2_keyboard,
      PS2_DAT_to_and_from_the_ps2_keyboard => PS2_DAT_to_and_from_the_ps2_keyboard,
      SPDIF_from_the_spu => SPDIF_from_the_spu,
      address_to_the_ext_flash => address_to_the_ext_flash,
      bidir_port_to_and_from_the_gpio0 => bidir_port_to_and_from_the_gpio0,
      data_to_and_from_the_ext_flash => data_to_and_from_the_ext_flash,
      out_port_from_the_led => out_port_from_the_led,
      out_port_from_the_led_7seg => out_port_from_the_led_7seg,
      read_n_to_the_ext_flash => read_n_to_the_ext_flash,
      rts_n_from_the_sysuart => rts_n_from_the_sysuart,
      select_n_to_the_ext_flash => select_n_to_the_ext_flash,
      txd_from_the_sysuart => txd_from_the_sysuart,
      video_bout_from_the_vga => video_bout_from_the_vga,
      video_enable_from_the_vga => video_enable_from_the_vga,
      video_gout_from_the_vga => video_gout_from_the_vga,
      video_hsync_n_from_the_vga => video_hsync_n_from_the_vga,
      video_rout_from_the_vga => video_rout_from_the_vga,
      video_vsync_n_from_the_vga => video_vsync_n_from_the_vga,
      write_n_to_the_ext_flash => write_n_to_the_ext_flash,
      zs_addr_from_the_sdram => zs_addr_from_the_sdram,
      zs_ba_from_the_sdram => zs_ba_from_the_sdram,
      zs_cas_n_from_the_sdram => zs_cas_n_from_the_sdram,
      zs_cke_from_the_sdram => zs_cke_from_the_sdram,
      zs_cs_n_from_the_sdram => zs_cs_n_from_the_sdram,
      zs_dq_to_and_from_the_sdram => zs_dq_to_and_from_the_sdram,
      zs_dqm_from_the_sdram => zs_dqm_from_the_sdram,
      zs_ras_n_from_the_sdram => zs_ras_n_from_the_sdram,
      zs_we_n_from_the_sdram => zs_we_n_from_the_sdram,
      MMC_CD_to_the_mmcdma => MMC_CD_to_the_mmcdma,
      MMC_SDI_to_the_mmcdma => MMC_SDI_to_the_mmcdma,
      MMC_WP_to_the_mmcdma => MMC_WP_to_the_mmcdma,
      clk_128fs_to_the_spu => clk_128fs_to_the_spu,
      core_clk => core_clk,
      cts_n_to_the_sysuart => cts_n_to_the_sysuart,
      in_port_to_the_dipsw => in_port_to_the_dipsw,
      in_port_to_the_psw => in_port_to_the_psw,
      peri_clk => peri_clk,
      reset_n => reset_n,
      rxd_to_the_sysuart => rxd_to_the_sysuart,
      video_clk_to_the_vga => video_clk_to_the_vga
    );


