��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނ�c���q�}�e>��%�(M�"�ު�hݬ��((ҩ�˻8��"BݐmV�Ӱ���dz�A�-��߫_�j��~	�Q&�Vi�V�V_�7�M�D��FL�?�q6���%�%�sC�8�㰂����r��l�+Ӫ��4_RR�G���VT���%����6���|�_��[���4&F���H�%Z��Y���qN��8<���mZ�{h(o�`]�UN�Yq��&V�Y~�ڔ�~�VK����7�* l��!�y������eKד�G�>�P��b��,�z�IV�hT�G2� U�� ki�OF�ނጕ�G�K$"ozr1Q^5H7�n�p���n����7� �mK�$���Tlj2�	�|$�
l{#�_ÜCt�FX�0	GD���;�@�p�N�VhF/\����l!���}��R��Xyk�8s)�v�F�3%��-t�d+�D��ApX�Kq�\���k|8��#%e�R�ӦY�CzR/�q��oE��H���FQ8L3�1ZS��K0���-�I�X0o=PA<��3r�X�ȹ-���0�a�5؅����j>W���IAu{��� ��2��Vt��4���.�,�\�6��<�?��%��ʣ	���0�Cr��]S��ʓ��C��H�<��S�����\yL]p�YN�!�b������@�I���;�/�f�Q^��Zޕ��H�}��!#*��x�Cde2�w��KE���S���7���Z� �}�k���±�gTV�̭�<@�=VG`Y+U���wM��%�C��!-��D���v"j�� "M����hDK�m�V�O�tz>�~����s�t��$*X!��ۧ�7�~oE��h14z7��n-������F���e�e^E�bP��2�I�ԓ<�:��n�N���Iݏt=`���nv&�K�7-�K�Qok�H�:ѯk��ĳj�N��s�2+�x�X,�U,=9ɔ��.��d�jX�-}����:k"��FG�&���J�mc��8L��W�.��(M�	���>H�%��w�%�߉�'v+&�Ťu�k�m�~9�=p1z.I�w�qC�mguao%-��������D��H,;i��(ؤ��z���v�u5y[n.���M���Y|8�&j��6��s���|�$�-ƺG�&�6�3.]��n-�͇�����?>��Ē.z��@x���n����ڽ`�[J��n>��/3j>�jK ?���T�yN �яNU&·�ؠ)�Y��W���q�ܓg���QvB��r-w�޲�CR���U����	q��+�=�DN���?���}���I7���6r����I���=��2M���u�A{��Sz�S�y�s ,J#'�b��
j?K�Os.n`�JP`Nz�>7.�5Bs�"��h�J:u�--�"禱=lk�Ѹn�(<��*��FO���ž+�Q�[�|?����\�S����{��+7��NW��8w�ʉz'L�<r��L����J�Y�DÄ��7r�a2!���(>�%�dC���f5)KgY�S�<��(����ޞ�]��i`��O}1c�d����v0���M�d�/�Ch��o��J��E)� ,��B?��F�����E5k��4`��3�,�*=����ر����L�3	t{kk��~y��%V�n�����Hh��h��_˹@�Sǒ��?��/�������kCI�)����c4�t���_�hNï�;m�`޶5�>;�B켾�o�rvh���x2�g���FK��f^�b"�G����צ\vF�Sg��B������2�C2�geː3����q_���w��������%��wo�9��9g�� �}f�n2�A�ޛ���v�#���-I l���R�ӟ؄%�3n	nY���F��̥�����)lq�g�a�i�_􎤓4�k����`?�vbu�Ҍ�X�
(���g��ъ~�� �>�T�G�N�*A{ΐ�]����h�`��#��K5�H�Ź�ɗ�2�������EĹ�X���W�~�]SH�6J� *�U\�y��g�8�����m�O��͖ל>2�{�G~t@-5�]��[�!1�={�w�<g��d�M��=�������b�_4r3��]"�b֎E���y�^vo��0;q�G���Z�7���dp�-[uQ�Oټi����4%K��!�S���� xi=~�
?�w �
H�$=GMΟ�jv�IЉ�?�t���O��U���n;$ɲԃ%}���]�RF��H�����x�9�I� ��pі�� #K8gm�Je�%�_��g(+\x{��窸\��0���/,>V�h��d��4e�� bfn�I�[D���X3�<R�D�P`^���� ��1����[�ҟo�
Ԉ���:�mā���%�M�:2+�:�W�QB��KD��(Lun���H��-��BM2j&3Q�.��1l�^WJ�P�c�&�?D�b/d�-G���kï��Y��5�@��5�5������=z���C �^αR�Ҹ4�g��9�g5�ۡ��E�U왶m~�p;�.�V���yR�Ƣ�T�y��\]�[E��ɇƱ;!Q����h'�$�ס<�qÐjuu���G���`����$�e�X���	^k[%�_C��h��<� ϧ=xݧ�����-C�L�^̨�C�\�<���^/E��;�c�~�_��jvֲ��;&*�]Lx��l$B�8��!�~	����K#��hOo!5���wZx�� @w!n1oy�ZV��<�;@�כ�OW5w�#]fE&e������`Z_���Sa{RU�4b�]������$J�R�<Z�治J��(�Kw^J&a����J�'�.Z�h��Ժ���K�(OrՖ�����i���Į����o���յ�����/5�M.ht�cƊ(�m��r�Yx�`b	��2O��(2�2�/bcQ4{#��k5Pu�)�o��O�E2+�1���4"��?ʨR;\��>o�R�o�	r��s��b-��p��QB��"� �3��Ŗ�C��{� p;��\����h��Vbꀣ��[����ͧ�W	�C����^6�C�G`�!B�y�E!.i�_Zc�*~�ET�׃%�����"&<~�!;�PY�~<3w�t�t�|$�<<E��<J��,K�aSG����� �q�^�qM���_J�9J�fɉ��^�S`p����<)�w�����^�7Q�ʾhQ*J\�EV1�B�Q6����<��D�Y��o2c�}C�Oi��-y{h���%�5ڍ��;\ �{(�12�Y�@�(�C֘�{��^�v��h���R����%� o��X._?>m�V&�'���g��"�n^ߗN6�$�ЇH.y��!J�����P�,����Mnt���EӞ��O^i����B�	��9�31�~�
E�,�B�x��I��q�$g���fkd�*���Ÿx��T�D{J�:�r���bhq��7�86Ƙ�o��cc'�\�
(��M�`�i��I�.�0���A`��w��R�T ��k�f�O4�$p��_ȉu#�`��P:Ifh�A��f�;X&,�a��
'�4�H��i�Eyr��(�s5~Zm��3'I�.-E��H9ǟ^H�v2􍂤���x�OV��ى'@���i��E�`�WH�'W=t����Q�a��Tj<
S�p��M�T��"o%3�i��AZ�d�+!8̳Qk�pr����4-�?O�^\�����	7!r8ddeN0u�ٌ�OZ�@g�x|r<5;�`�����}1Y��	�9��A<��R�_��e@{p��el���T7�h�F��@�f�s��SG��� ���m7Y�����-�l��3Yb<���0�A�ý��I;#�Ev����u^�rLk�~�����JI��쟧���N	5�9��0k�� /9԰(����i��h����i�-�� ��A�G���y7�\z�l��`�.Kr�v�U��<сEz�noyhz;\���B�o��Nۨ��L��X?�����;};�e���*������3��b�4Z.��9]Ä=,V۔��Gqx��-��e�ѰWo�ozi��q��(tS�J07��X�X�d�=I�.`�J��w\��4߷��tT�D?���U(���L�+��@�Ɓ���Ѹ}�1��5����&��Dò}��r`�2���vb�~΍�І�h�C�o�$�5�r�]�GN-=7c�W�ʨ�]k��Y�_�^�ζ�'P'|�����ȣa�s�P�vf��-Ƴ��h�vo-����z��).���؜�H�,��RWq��H�j�V�P�H��/�}M��X������|�iJ�L�<] ��Z��1*�P��c-�-��:�q%��`�ݭ���t�;������-fL�*	�Da+^�%ٹ\��a{�0��8����J���!H_f�
�i���==�g����/��:!Z޸�^����ޞW�e�i���5!��ݜ�,z�f��4-�����n�]���l^���~�~�P���L�kCV/+���wF<2&ל�bq4��s�L�<$aH=�`��}2~�6n�	���,k��S�Hⵎ��N! Q��a@��L�[��V��'6��-�� ˧�X��*��ԢWPy^٧""�j�)Aq���94��:g�R-�D�|�-���Ɏ�7�\{�۳&�~z�i0�����M���sk�bA�s����|`���ΐlWk��C�����U�_�Q/�$K k�C=���I^ͦ���
yl:�R9B�ĉ61o7#��V��v����˓���r��IH'~B%�Y*��yx^�M�౬ҍ�[��U9[#u���0�V��Q@[�c�x�#"ލIT��-�x�+���.(/8jዒ�y��'�Q�!�R2����J�-� �72��e_�ӳ�pЂ�!�\�]`{�8n�k6�?�������Ţ��)�O&�R�\%�p׽��]�+�}�c����Չ��x'���~wd�D2�-�\��KT���n�0j�)�/`�c���I�ԫ�X��u\����m�RUno��lu;zv%zRc��f~t+�b΂\0�?��>�<)�w�8S=LXP����Ζ��5�%�5��(�`����zс�8�Vj5��n#���9l��0������Y���"̈�P�ٮ?i����'?�W5��L2�*��°���;�-ӯ%���I�5�w�t�\�򙿲h`D\�C��"��L��ɦ>��]�5��w�zZ���&r�����Q��I˴Z\p�����i����2���f�|�d����@D\�ֆj��zs�+���'�7ϯ�2V�Z<���._-�����Ⱦ`xE5�Dt�T�ĉH�Rz��`b��҇hv��F?�8(���Wפ�;����r>���M��� �,�/�D���색bDp4���J�ag|�w.�2D���3���S��
�H�~�千]d� ��M�p�N�S��)w�^���'�f��k�o̐��8���&��^��|�k���O�>J5���{�U^��(!*f]` UP�W��u�| .{f�j��xIUL��q�&&/B&5@S����M�9
�u��ݐ<���#�D��|=Ѕ$ �� �`�pzD�J4���f�j͂���n�lc�������/Z���S�|�*D��S�jw�\��Zw�5�W*�37f���P.Z!��*����i�2��;ܓ+��<1���Cf逤�֏͡R"��U�0�Ar��T4'�ͨ�-?du���*�4dA!&�̜:F��vJy��w���{i�Z��K5�Iv(�4Zjѕ�3]{ˢ��Db�;�׍���ƻ�B3&z��P�c�'3�� d(ZQ�=��[�2;^�ӕŪ�J�\��Uw)�za;��"��GSKҀj[���M�0ν�9�A�� D�ON
s�T�/i�Y��d�'�nL�
�PW	n�����,�Ʒ<1)����O9Z��eoE̯�J�ߵ�Ǿ�C^����p�PRZ>}���g20rY�ܢ0�n��Mqi7�k݃�jf×~>͘,}W[��Y'bP���٪���ڗ���s��K��UC#䫘_vo�9Ct�l�|��Xe ����,t
H�j�����5��+))��10�� R̍[�8�#�,w�g���=W��1�E��A�T�%ze@���\��Ux�bZ��K�p��i>�����жL�J*;pc�l��cQS���J��Q�o�=g7�D�틇�\������dX_��યD���1a�yH����Ј�D�`���~�T{H�6`�]3^T^��rj>o��Wo����`,�⡮ KK7�;n�3�説�h}��Ta�dQe���4qY+��=�{.!��N��)F��~ݒ�T�97ͪǥ�ִ��6.�s�./��#�Kcy���2d�gu_B&����;G��d�釗� bƔ]�cO3�Z��L}⪗���2L,�L*g��O�ܭnm$�P\�Lzs��������އ��9M˾��7̿���T����|��)��ij3��ȩi	���S�������u�v;LP��. <����Yؓ[��W�ۙ���:B/�\zl}C�x���	�,VX -� 0��;�euŹ�����5i����0C��լ���.��]Y���m�?��4��N�R'|]R�=K:OMZ��"_�i�]�`�������P�"��o�?��âi1c��yhl~Ԝ�P&mK���\պ�Z�Cͽ���4잤X��I�t�R""�8�g[[L��Y>�T��HuD���_�dx"ȇ��)���2����O(���t�m,�7�HL�J��e1�ȉy�n�o/�:˖�٧2'�L���մ���j��U�PT\�4�|�I4�����'2��y\{F��z�rw}�T���Zգ��(���gz<-q�`�ҿ��<��,��;��9 �?
t.�c�J�d�[�R����+���V�9���R�j}�R+s��ޒj�r��9{���z'�8--��W�b-����������0�s�F&��� �Iw����GAO�鍰n�i	����sA�_5Q������$����E��Ŷ���K�B��	��S.�'��I-$��"���_.���:U����[�F��D�6	������Z���Ƌ}j�C�@�ޠEYx�k��qk���>L bR�+�
U[�36O�B�fxХ��qZ�Hg���ب��4j;3�O��mP�J�D���߳y�P�
���*'�==�8�����)x6�¥&fj����a�<� Zwݣ���ܱ�[����:���޺/%���2��<�#]��$�ƣ �	eءZ���Dar�:��!^���;�`
�������k��C8�te;>?'U��K��M�}�mѫ��X5w>)������k�1-��d��׬�^l���i�W���bU���y�0f(��T㟎Ъ �HM@]m���"���%��!�W��~�K��j����1����rG2$����3�f	r;P;�*[6D�ݮ���D3{_�%xN�!�s��0Yo��a�u�$�ņw@�(�k�=�c��w$�̎���ۓ`[�>�����2z�_�n����їIGb��
�n�����a7��v��>"�N��γ�9�3�5VOKo�6�
G�oX#[��!s��Q�P��#�]ұy�2o����
�4]w%�r�
=�5�0��V�2������2Č2W�u�9]�����V�EΝyO��L��m�H]�ف��g��N���{4΃uj��&J,"�T��$'Q��͹'�:x�6�3ѽ��L+�c��rQ�J����a���`��ut�c�F��T[��a���#4xO��a��Ԗ�f��;����m1��Zb�͌����S��
�+ą����;��ezW3�q���|K�I*u)k5�2����Ĕ������77��0!F���
�ZȌ��v�f�=.9�`��z��&K�tM�~φv��E&����k�᳭�]6����+�@٭	�9�/�5hl��w��������Q��2~i��J�yo��_���� ��yv̒������cuw�ƣQ�+��2���e1'�	��L����y�0p^ ������{����x�,"ΐQ+٘���w�d�#�g��q�l���i��c��x�̚�uQ�m䆂�{��/�����KD������R]�ҜK;�14���������Z�w�g��i&�o��n+��%kC������_�ɲ�,;{#[�egZ`�m�y؁�B�ڴRB�i+���с�.V���"���r�2yC�c?^�8�y*qP�"D@�.��RA���/95P	QWfb���v�z@O��ϚtYgi��p%߀w�6�J�GM��WHrU�o˖��g�.癨���&����`�1�mT�B��a�"�~���7��2�B�W�����㎷�ӕ*{�9��Zd՞�?�w�b]&IKtڸ��y�i��>�#^.b�=Æb"� �O�I� l���<�D���vc�(1���x�b		Y��=_��B{����C��Ζ38�ʙ(-+Z���/�Y���wp�8�?�\���3Ϫ�'�n���Y7��'e�i�>rV"�q�l �RTGk�jz�>���V�3��;�%]��lx�N3�?<�@�>�tj>C�|YOZb��ןEFv�9fF���l�L�t��SR�jО�^�%ktw�0㮩�Fc�0���$�a.luk�2Җ)3����{m��	����?���<-)���ɏ��
]8����O�%9��2�PlIa�$�]ק�썇x����~� ��/���(A��N���Ž�hx������d�:�bk97]�h�?�9 �<i.qCE�sy����Ń�J�lC��ڜ���ɺ�=���7�|D�}0�s��D�\��q�1�@o�/x�� u:��D��:7 |�,�	�k��$��{��6���0�n�N���JA̑ğ���=�,�����?�.5��,$Q�͔�!�:�z����H��H��Fi���~��b	��#L�[,%|�����q��j�f�$�ߣ���uY��#,u�q�m���K(t�hnֻ&�ګ^��[����DT�|�U����/����:r���K��6`"���z���*n|�m�
��¦f�`�f]X�ި�^z��
O=�gB������j3�^qI�O�?j��.��}�5}!K/E�5b�P*�l�Rn*Ś�eY[��&�!�%��J��B��!|�5���fE,�Ͽ�� �1��Ɠ�b�썔�\m�I}.���)��:p��hˆ'��L�&A�̾�)j	���st������&���*q��O���U&�L��m�	?!�1��W�H�S�!�t�9Za�mC�G�x�A(�,]��_GdD�钛�2�_z\�ʉ��%dSXS!+��2����Pt&<��B�|.06%LIR�������K?MA�$��n�Կ�����\#c_I��<�qw�I!`@)cB�Fr�8!kM�
�5�i�^9=N`;
S�ةr��cw�m׸<<�Y��%�P_poG�UŌ���4��W�5���eԫ��%	̉���sl�P!wđ� D�å��6�Z������"��ԟ�Ϙy�!���q
�N�J�Tx�P�v^ﺖt�K%�<F�
�e��TK���'���Lp1B�џ�|�� ��! �޵%U�c����5�E*���I����-�έpڷ#�$buȓd�.��H��4h�y��IU�.=:�(�4D�biTb��~�m���k����^��T*0x��Npo��b��� �F��<��Q��o?�S�������Q�	Q}Ւ��)5@q�ZI�n�eJ��SrD����H74��`
 <���WFm�aTa$���!��'�`��1��8��05�2a8o:�^��w����s������;�`�h�������"�]"N�Drj^|�fͻ`����J�9,V�QG������xG�� j�oc�E�Q�� ]_3��Y�
�Q���(�U����8N�5�����$�[ ��9�1ғƧR*��)p��E\4�h�P�Y&�]���4E�}�+ٍ�F����w!�S(n��C����`R�����Ȍ8��.�/������d�[�mf�Fj��V�ӭ�	RŦRQ7�Y9DN���-��y��P��	A��+n��'r�O�=���� �e�	�"�
u0����ȼ���Va��s����G:Rҩ v�h,af�r�e�F�͍e�NȌ�EU��2'�������h��;u"�F���ɓ�B�	ܔ��:6�"���zh��"4�i�reK~6o9��v$� �S�Sx��u
t]E�\��x��F�����\�'ي��`1~���+�l���"!����M*}W�:�A�!���9I�Y�[��:|rD	=�bK�������І e��L�� �}� ���DK����s;,�LZ�����C�����<��	,�%�k��fn�Z��?�ޗ�M���V��
*B��T
-{�h��z@�W<���׳�!�+Y���9�X<졒���0t���ם&�Z<Gz��W���ڟ-_�i������}/����#8��v�m��W.R�2��g�����)�J�Be�s+�ᰭ����[^����a�Y�L��~�)WwU��`1���ID��s_ �ϲ�Λ�2l
]u�������>��Z��H�]�g=�dZkE���{�t�K0�oܽ��K� �r�⎰�7+�[@X7��;�7���^�{���y]n��}�u6�5*+̗C�ݥաC�[�n�Aa����l5�T�K�����"�p<EC4;[m�+)dv!�ȁ�f�̍�FjR��9J24>�l���w�ֱ^$����h���5
�"Xx�h���\F��jgӾ�'� H�����L	�'c����G�\��A���K�D��1{JxlU��9�P_�Od����dΤ��]�k�w
��š	�������f����K:
hq�E��Q��|([9���0	�O�A�s�F�if� ��3Ӭ|E'��g�Sͷψ$@B\�\��G��ӡ�ר�#��R8�/�5�e��q�2+�.�u�P$@u-�Xb��U�4�{?�I�,	� ��=x�_��q�s2�J���M6F��AT�Ml)G�m���]���Q�⿩]}��,\0��Csr���i��q�9�cw
6�b|��(��E���*�?��;^F�A�y��;�h��ݬ��:/ivA���4
P^n>����y��~���~-�o����&ר���(C8k��v�<��դ֨K��Z`�#K�\R���Ά��m���lP��$��R!xI�e�a7E����)J���I����o�6�IC��0��f6�H� �WW��4�"!j�軲���� �`<�i�+��
9���uzg�>����/�+��|,J��X�w���xkd�N�k��:�Z�Yz���{��,�;��Ʃ'�z���#�*e�%)�RM3��SI��Ւ�8��q��_�{d"��a������QFk�o٨��w���!�b�MsG��m��gͻIi�!c@G�"��c� L�X½�䜨�@��O�v��c�)�7���d&B%o������usA��0�(�(����>_�����f�"���(����L��Gd��J���ʓ� ~�/W�����b�>4EnGY1�!PUV	.9L�~=��9C��N�]���d	�S��
���V�`S������!#�RW�/�A�Ah�7�u@�z�T��`'�/���9ݍ�(/+�W)�`3�͐^�NƜ&jnZM�w[|h6����z��i�i�_3���9����%e��8~�X���F��Ik5������p�̄`���a��o6�(.z4�A
P$�i'�?�,�����������Ն{ے�6�_1��vXԨl��O�G=�r������}T�6k�Wڀף�F�	�j��o���h5mcVMd��Bf@$�>���ڬ���൥�WD::�����C�s�����o�< ,��X����$˟-����4�r�׫�n�`����h03�;9i$��]��*�<!ٺ����#������ʌy]NK�!���e?���]k;��\B����s^��x�"��ߵs��{�놟�Yщ�\\��71D%��%�N�]s���Q��(+��蠌b�眡����Lg�y�FPJњ
S��\��9]�`�Q>&L(�j7�t���?t:rK����h���s�#B��r�'���ll�#�Ӱ�/bт��4�}\މ;syb������3U�2��e�P�E��s��67� #|&(cS ����ξ� XJ}�`��p_��M N����H���Ud^*DwƑ��+(޲<�L�S'��x5_-;Z��L��T���c{��կ�����]�6�.�+0�|��S��\+puiN��+ф%^����"��$&"��Ӎ���dsγڥ���L���_{��f.+�|!�����Wf�	b4��_F�0t�l�W���/�n�����k�P��L.[�������ǥ�
��\��s�C�fj��L	��M�2��GGg�m�7�[���J+`����(�	��d�L��v�SM ���Z�_ْ��BI,:��H�V��ommɩ��u@3�+L�Au�Qŏ�ԥ�ui)�yZ,��Sf��
�<a�M�c;.�����<g#=12�]Cq����*�z�N/��D����m#�T�<+���,�	l�U� v,�iMd�ݬV �%��8��Y�bY�h`a@%����'X[`�WI�G߸�u�n�
#���F-��ޤ�Ő�mW��!��Fù�����q���w�-�=�}	iyz�*v����ݙ��k	�5S80O�/}�j��������>�g�S��^^8�Z}.�NR����V@
������f8s���^#ޏ9��\B���>���{i��t:Hx`�v8�{�e'��և�I�,�P4�����]Q�w� ���;�^��MR8�GVt���2�]�`�R���B��o��7Y=��e�_S��F^{턡C�L�~�3h8
��G6���#$���[`4"�~%#ʫ��p|�U��N�GӪ�o��5��}��wd)X���B�UB�_����×"�
�Y7.��yta��d��6[�f%����%�x�X�Q#p,�O�A������,��,D��2vm����Ur4�G�
u{Bת����%)����w����CZ�;K� �����=ި��3<�t1����-8�&Pw��<2d��� {!
�v�×��#Z-��U�X̦/��_��=���EO���W�20��pb�6?��)X�lE�I.�����&6�1�C)����{D�U���1X���1�c`Р*�4nf���芿^��gB �D��%��� ��r��'�Я���B#��!�"Y��>�k>���̍g��c0N�2dM���䝔��#���T��Z�w:��7��&ނ�mut�c�ңd�ξ�e+,��h��5�J4��O�$���Prq�_߼.K���5&Ch��&����Tt;�:H��0Tc�N��Ba��d?e�_�8W�_9���i4p^�j.)����^�aBc�Kr�s��%�^x7|��f�����
y����6Z�������8Y{r�{!E�ND���v�"�D�{��6cϘ�S(��)V��h�80�5U�µ�J9�[|M�U�e��m1�.�t7�]�f�Gu+�"$��_#]���^�K��f[�_e��0+.l�|��9�ɾb���u��6���D�IN��;��Gk�<f���5`���O�F(	�0V������B,��u��5+�Y���E��ZovDSgm���t��#v:�ϐ�v(:4�	�]a�E -�mg-V3M[�0����7�F��_I�8E����05�io4��<eU�������H���6�,oKjr��G�.m�B�B��w�&�Uu1�U�6.����������bŰ �1�z
v+6�}�L��=1ќ���/(8	G��=���7Z�*Y�7No$�m���&~F��͈���`��m�V�U �`��s�Y�:6-n������e��H�{�vGS�0��֪����vQ6'�H�6{)����X�fr�r��%�y��L?*;��o��>2>m��ِ��������]z�| ����co*���K��s�:���A�0r�4����
s����pU���<�o���B���\���7d���N6R�k�Fn*�9����k�@�vk��Jqe@ų{��d�"k#o�ٗ��J��-���OX{Z�B��c2V���˅�G�#��m��N��eT6ɧx���6�[��q�n���<�(q#����������Gf~�U�u�`��}�G��T������r��$���N ��̐�u+�A��pH)<��j�jݚ�Q���&�K��N�Tx�[͋�Pc�H���چ�'�xUȫ�:�c�u`Z�ج� �,�v�c,�!�ĸ���?�i�;�{�ہ�Q�aN��O���j�J��Bp���E�`(N-g�0w*�yVy��I�BjX�N�E9.��w�X�TW�ߘ�;���|g:������/�Mmp�"	rMYX�╫����G�;$��A8M(�������=y$m4��-YɸñV&�"	����O%eLS'"ő<��>�&&���"$��|�?�f��J��� Ч鐃C߂;ЮA������F�8��c�	c;�M⦣�A����!���,,B�l�a���#`]�v2G�-�4�Y]��<�%��ٴ�8��
@:�=�m/T��ܠ*J��vʱ�.�uU���_U݄���<V��n|~���^�]D��x���A�P5����o z��=���9j�>�O�H��m��<>��h���dv`�/)%dJf����vν3$t�*�c�r�����k/��J���k|f�V�*�HW�;�5�%�I��-��v/�2�ZK�vW@�L��U�(���,���17V��gS�X�D-}���yS) �  g����],$��Kl����iQ�9^�)!�%;��_��1���2�"u��kL}=���	vص��>s=���E�Nb��.��A�k�~ҝ��m��_�%��U�%!h�5�d�_��%��r���s��P�<@R�t%�6�6V�EYv����=�����&��8ki�F�i��㻮������$�~z걁��y��b,���OT�������H�2JH���g�羺*�_��/A]@�~�3Az���K��(�_.?JECL�{۸!�{6��/p�?�]Q w�@���M��`�{�V�]T�v�	��bc�����V�32��_É�.E��0кT��˘�k=�C���il[pk� �LK0:��=���z>пU�d�������Sc-eQ��;����Kv
�6ea	:��$B)íe5A{C7J= ��ha\��"��1I5����]��钍n��)��!>SOX�q��w(~��p�F{f�wh�\J��r��fs{��aE�۫E�@J�y��G� 5����~�%��M:a�-y�I�jWT�C�	����cc��n+��^�5'q��i�3U�}�� ��h���Q0���m��`��b9�/��C N�	;Z�r;&����/�-�5�5���ұ~��Y5ih�z�0��>m�,l�O/}M\w:�By�kfP�Y��H�n����u\pr��]rtD�����$�Ԉs�:zT�ʯ*�zU4�֧����n��s���
s����Z�Ix���D�֚c�צ�U�g�t��=��\�;{�����1`����s�/~	��Q�q�݉_�3oV+I�����G�ԃo���������}�}c�nq�. \X��0�薚��S"d)�ć�+u�P/�NW�9�E.��6���B�<QE����Ǣ��:�
\�"����~�"�x\��ܖl� ���y����j���1`j�=�(�&m�j�>n:ФV%%|ǰ����cE�� ST�|CrjQ����]���zL����Q�`9������d<]���;�S=c�%��Kg�U;F8K����?�^3%��2��̗�*�5�@�T3k
NL�C/k�s�d�x��7��a��gXu��;E���xù��%��E�t���B=�:3��v$C7���]��I2�`��Q��A.�ڬ����3.,�8����-�mSw�ŹL�q@-aB7���k��� ���{��[7�f�$�*D�rV�����)�:9���u�}��.X�F��mn�R��-1���Z�&iE\` 'B����\M �5	�';��6i;���H�9oXBN��_���3�q�a�7�-��I�/(�[�;�y:>]-(n�vE�Y�_��3���@UT��>���jsQ��F�#5D-�>�D��*8���b��' C����Č�-㤓����4ف�$��@��T�Q�e�8�E�#7����n��<S|�aGy�&|:�xG���u��Hh����#-H��1�0~��qe6/�wz�r������WR����3|E?�����������L��'��ga��l��gAj��)Ӄ�NlY�c���ꔴ��DU�Ĺoa+�0�wA���MV��������<[O}���$��T_��(��X��cﳱ��H��Z�����c����K@����[��ܶ(�د����d9r1g~�C�����e<)�r���F�ڪH�N�=�p6:�I�l݉@��&PMF�v�J������{ɽ�������Lw��P21�\��vYMM�0:��4k���s���Mf��a���J��"sdT�K.������u��K���oNݰ���kB)`dc���
�)��1�	?�nȥ]��I��,��\��� y�N��%5���1K/��q�e�}+��N|��z�R��67e"4����%~t�W� B+rY�a$x�{���~���/ 7<�1�[ę��'�W���|�&X8��]�*�ǝ�g�n'+Ln�E�ˡ�#�g�g�x_�;�n�����e��o�W�R��sp�R��W6S)�G�ڼ�m��/�eo�_z��7�J�����=�iݽ?��\�U�������}.��/��#����
���꧗"7n�*R�	A���M�FG+=t�>�Fd�b�8��T٣�MO3���~�c�8M�z��Uh'7fr��s��	�-�E-3��|}'�o�So�:���������g�[Wa�AI�2ËsL&4��
�u�}�{~K�`����>�~�7C�xW5��wm�c�ꉣZ�1K��N{2��\m�R��(�t����W����g���/��z��ԐMA��װVd�e�ۑ<��z��D��,�Qj�k`�C�^���FY*��M�P��N.�?ſ->r�]T�+)�xDT�Y�y|
%�c�͋a+@'NX��Jt_���Nkϫ'��2�%��/b�/��E��;V��{��b5VrbD���0jQ?P��M5�m���N��d�3��+�݃8�9}�.�F0�Q�pQ����]����yG�3���9�?��d�0j
p�v�O��[Q���<��6�[���gO��������𡝸۝Z�6�s���p�d�����M7ctT�YP�̡�S�#��G�U�?�8���z��Щ��ӓ�/?t:�+��μV�3Ꙛf�J�L8Vp���uo�wę��	�fw���o0S[FT�B���m��r9i��#u�酴�g4X���*1���A����͕o��~�E���ΚZ��I�q+BI'���1�cQȃ~� ]S�\o�7-��-GQ����M�X������C���ߝ�n�r,:�U�^p0'3	r.�M&�~O��'��R*�}�S��A��B�0��M�����E)uWQ�d!]6�C�n6,H��F�O�����^���
��[��Y �R�gk0;��*�e��a�a�WA�4�h}՜�y��?~�E�:Qf��e������k�̩�C�|
��D�ד�`��Y\YGSe=y�ώH`gDQB�l����@�P`<�P���~�G�&G�C�L�X���-�G;�J��5	ׂ^A`������x�;Y� �q3�p��`k�ٜuu�NY�[X`Os��5��.kt�,�M�VvK�-��Np`�Io�ov�1[ϝ�I�s$DD��BS�s�(��'�s���ټs�R$�jO&\�@���v�R���a��>F��� R���j����|JH-u���yA\'|���/*��k|UW{t�[D�R�G��^�7�61���?e�8�U�ܯ�M��J�#A�-t�x/nz���Z�=S�<�\~����:5���_��|R=��q���������3h�����.t�.JR�қK�w��[�WA�?�~�qx�bh��"B��;ٻ�b��X�zp��ݶU����t�K.��)<@W�k�.�۔�/�����D��@�+�A�d���я�34`����!��_���zX$�f���Mӵ�������6���v�����:��d�������T���9&��Ι��	
�g��;%��M���Ǝ���}�/E���@�m��Ɣi5�To�/���e�[�9yk78|�Cy�Z��UT�H�\5/܏L�6-�L6��5�Ϳt��&��5
��E�ĄG8�eC�j�x��_Th�L��A��S�?��JU����q���=f�o��>��,/�=�� ?��_���=���@ĪNT�K`ɣ
�e�/q�g��u:zDn2�A����ژ�jK^8��w�H�/��-|�B�7��[�n��}DD�YlĬ�+�{�DX;��*z�49���-�D�R��1��V��Qy���/m2�)D�qD�cv6}{��rjHw��&�� ���+���_˫Qߠ)z��>L�C�L�(�V��l˝�����N��܄��<'�EX�a�}�p�����@��-Ȼt�ց|�w����#��gV�wn/��:R�2��������hv�4��`Mo��р�H`��W��|���RtO��V�W&il����~?���]N�#�g���C]��<���[.�0]�W3��د����q�\[-.(�=I�}�9 ���ŀb�W�1OߑrlQL�4~�c�Wn��21~�`=�|ũ"�yz��rU���qZSVo���Kڼ$�%R�U6���l5�F�S�8���O�"O`^�y��1(�;�K��O!�Ū�;Gis@z-�h�2h�w��W^ �����J���F[F0�g��>�,�x��_4%�3�˄�Ir�c_���B�5[RO0�)h?�W��ڪg�m��Ύ���JOfl|TW�&J��I,!�_ʣ��2�״ԟTQ�}��Se6��1},y���I?�\H���͇C��U���l#���Ό�Ɍ9".%il\��<��-F�Aߖf�1 ����A��4zA���POK�Y-$�G)����j���_d��� �����V��_�&�1�A����^a����5U�闩�87����򏦪��	�?a@XХB,#���ZL�r��L�3ll�p�6P�q���n�=fK�ܚH���lX�� 5�A���7��i3)��u�oG����,gT�ح!�#s��5-'����W.-�f����3������e�����R��4�5׼z��Y�il�3���'h�E��]��	��Y@����=~�0�X���*�E뒱*w�]y�����{� ���|��D_O@�T;��L�����z�O{������Mjq�ʰ�R�e���B�Q�d <��Q���A���2Z�-��o5o&(ly�tx��ȾI	�D^�����Bu� �/D��g$���$`���6�/����VHPww�=u��cA:>�T��X��P���dF7�ڄ~���-o�����:��l+���!��/}�jX}f����u�R��}���dޝ'���i����W�;�s��,�]��ү��y�[��}q�a��GW,�'�~�e�s5�(�-�|}���-�O�;۱�>�;�0��W�_'VQ�b���"�T鹋~��T�kF4����^m�G|��"�\�%F�=��xW��\�]��v�,ܬx0e�Z�W�A����	���E�
��_��OZ��h9�V\^I�Kc�Yr/�[�*;�`(t�.�8kȾ�{�e61�ٛN��ِQ~�`D�#���[�����Ż�gk�\�.�e\P�)���)r�K��41���b�_�T[.�\�z�R��L�H��P3X-r#2�>�*z]69S�W���� �M� ��u^�%�����m� �g�)\X�!���/p���(@�4���3�T��i���	�M����㒻�V��ܢ`%*<%��i�o������¹)z�o�ϱ(���:��e�S#��%���EX�*�tp����?�<�Og�I�m��^�c�kiV�:��Ȝ�u���ei���0�����5�;�jv_�Ďm�?��$��I���ΰ2�(����=yg�g�>��d��BF��[�{.�6���lm4���F�K��uh���������
%Ad��ʆ�G����h�Xm_ri�G�GI�CYAk���� 3�r]��RV�]��7M���wlR��BI8�	8�K;+U�ӑ�go�ma��No����<��w��^�(�����^4*M���Z����vf�E�
VJ6��Vp���s��\"zn�����BW����iE�V:��^5
��Z��	u��H��\��W�4�no���� �D���o2ĦF� �G.��F[��0�)���|�q:>���,k��;x�_�DiK�2�QW^O.����5�@@�Y0�=�H��|P�S�WD,����G�ݛji��b7��]������K���6{k����Pq{q!#�Zk�?w���b�7k-�o)��C;=���S!Q�q���*Ó�N����c=��֍ֺ�E?�h{Đ�f�/�sMj��R��a��g���� ?�¢#f
Y�%[��̔�n��`���W[�ȯ�)�\t4���54O׆�����h�}���ʚt�x���ig=�T��

6b]��h�N-�Lj�[a����?�{)r�jʡCg���j��mp˵�e�#�Ua�R�O d�fo�ڥ��h;&�8v�,�hv؉��jӔ��ZK����T��j�$e���ڶN�!�ޑn�� 7�������UW �M]�d�Ҽ���]51p�#}�z�"��������x�I�C�f�Ss��&�|R��!J���%9i��(�U�^݄;��+���)_%���6���|�m ��x�@�E6٠�*7�N��:��{��� �P��YJ�?�*��J?���YZJ�����|���p�	J,�h�MտW#_M	�X�>�"8{ÓV���>lY�����l��� ����G�ߩU\m+2-ǋ�$g@�f�^�f�ImӅ�B����r�ſ�]��`(��	_�����%$��^W�X+��7�H�?�oPb]}>E�ᠫ�A�EQ�7��s�g7ك�X����D)�}�ޟ�	��� z�j�Ph֔���x��=�S����<]vLs��L7��(u�z���&^;����v'9���W�a�K�:]ΐ�.�
B�
�v�����1�;n�
���8�jh�����(�0�~H.��P&|�1y�Ao��9��A�U��H�g��b�9�}�7l��+W� wӺʨ|K����x_u�O�b�� &q�>@�T����;�b��_!��C3`���h*9���?Z8s�4r{!���&�ƪ���7�O!�M����yl���ů����M�)�V�>��:F�`���Ǉ�}Qٻo��gog�?PV]C����1>���&�q<��"m�ƥe�r����ǒF@��]7㕊`E$�I��E[1��k�з&�!�ܴ�N���Ju��t@�ƌ�C�r���`\a� �C�[�S�i8������R^���;�� ���,�:�ӕ�#���v=�ÿ�5.����l���{{�g���A&������_&�������e.�h��f�5�9�&�a��=Y�߼V� HE�L��ژ����#�$���
�z(�o��hr�l)Y�XZ\ZD�9g��x/�S(iu�����/����+��\S������%~[�*V�lc�C�(9�Kʒ�� ܪ$�Ry]&/���(-����<qu�5��_7�?�sW�H���;h-nCyO�(%����{P���Md��eA��F�MWR9���]��J��g�r�f���U}v�~
g��:�M�YY7"P�<��6\'�M���,�p�I�ۭtl�ȑ�dJ�s��*Z�C�9�C�ǿh�ѳx]VO[��9��5V.'�
3 ��!����-B�8�u��{Ɨ���`��S�1p���!fyP0�"��$Q2�$�2q<��K}�aH��ߩ}�I��u��YO9�.����w��DZ�R��庞�.����\9-e�-�����!Y3��a0�<��=>����J��HL����&"&�ϐ��Q^��	~�Lu��<�L�M�� &jo%�Q�$ٕ�[l*��;��+�_��z;�t�?�z	�'�c�0^�p�|H	��6�����Ed���!���$6wcZ��[��5����_�Ӵ�'c��
�c��`{Wt��棱X
u��Ugsc��������.�%�_�0�u9�W<�1g���7Q0�/�c�/u�u��Ɲ��f������3�� %}�>�	�6��n�����ǟ`�8٠���"Ve�k�夬v�����^I�A��YAӷ��3�����ˬ}�W#G!E+l�U)���O�O�D�,���B!��zD�q+t�hw�|h�JʽR�iU˚�R�O-s�q`鄠�M��ıVd��x̑��%�]ߙ��w����BA����C5l:1� �&���h�r���	AC��F�����	
��: ���S�+V���_�p$���h���:����W�@�ǈW��.�����P���S������5%E�h��:b^�|M**��b��J��/,hl{j<�S�ݛ��b��/�0��Z�w۶��h���C0�V6r4��f_�d <��6�7�,��P�}�u#m$2-i@� :JZ���VF�/G�m{�6W-�-8u%g/�l��ZSk7.�X���YVa-���Szo��9T-
kC�_��Nv��RNf�R8K��$~��6��'G�rKȍ��ރ�ު>G�꒣K걪)�������V��Ӊ?�(�t{�`x�զ�	0ޜ��p>~BS�'u@�a���-�ܔ�:p�1�F����V�#:�����~��Q��X�����sa��TJgd��V5����	���[�����������7a�:߆r�i	�YX���/�pT��7�!%oGݑ�p���K�m�;'k�B�~�z���o&W�S}RT�����_��B���zͶF3I�~��(��z�F'�S���$��@��z���w}I��&���c�l�"����+j�Y������b��c���W����Ij���S)	�l�M�wF��R2/E�Qx�0U��˾��r�`]�ֿ��Ѥ�B�����W���D~Іr9�o���//�»~��~(D�����e��M���:��+*?��)�濊��Cp;�6r�
;2�8M�^7 Y�E��y"c_���s�r���U@�.��1/秶^`���y�<}���p�IJ§��j�Oi�me�Xp�����KE�3w�K�!�-�vջ"@�B����/���F?�□�T���1��RLy^ˊ<�`e)���0���� �`�N���
�����TrB�q������ G�ڒ�������U��dR�*彖e�4�XU�1��=��4w��P��	��2#<y��Mn���O��&ߊiȃ�F��*^Uմ)C��'����M�lFtр�zj��.�վM�vv�d1A�q���.�����s��No��,�iw�����o�(+tQ�(�p[�G%��	�"�L)�����J.q���s;��L��zX�kcr�ܼ3@0�}�8%���!�9P4����b`u4B�(��q�	�A�N��wlφ�P]|��e��c�Sy�)Z�V*O]j��/Q��Lp��SF.�����E"<��1%԰S�@���_�]�];{ѽ꽖�%�ZolD�v�\���i��O{�Q�E`����R��ɻlL�r�?W�NF�$��x�����kվ�W�@�wg�W�d�38��юF�e�[K߁���~5�����
I>����)k�s�m��Ȓ.O�)6�SݞtšX��1(��L-��ϖiH=�f��_J��4������f�{SE�Qp�Ѩ;'y1�d�h��W���Mj,uԑ�h���6���ҽ%�!���5.����~����OY�XP�v-g��E�EQx���r�wMߢ�f���S&��۟p��f�xE��3u*A��I0�����N�B��}���Zᮼ��eGrUb�8f�j�p9w�c���{T+~�U��[���ǒ1V��OB]$�`�WT5�h���:=�̃Ҧ���D㫱�ѾZ���&/�v��J���J>ͯH[��c���B���+Kx���{[o�MJ��¿�2u�.p�#ۻ��"9��*�i}�DF�=�'Ea�ތ㇕�{�Н/�9�gpH}d?�(�������
��}>���]6PM6�O�x�hzJI��|&��S�L���ч�4�7�D��S�Xz9�Yu���#g�lV[��5o��I#@DѮ��qsw%E�z-��x�����s��&���T�J*�܆�#[J⥃���%����,����h/���jxw�Bn5��gu����k5��A�����,�m�M1�r��B^��"��19e�_��۝&�eu�Fw#�l0�"���BJ��Τs��l5U������J�Z3u�'n�\_�*�әƈ��ӹ�^�-��V����f-���U׭F�� ��F�ms��A�QG����ҫ�Z�}� �d��|�(v�(�����|9�J�R@��^�y� �#��S�v�O��~&ի� mA2��� �YҚ.&�>����to�����Qm)�+��l��wl{�%�^<��3�-��t�7dY�a�J-z�e�Q��iӳ�����`���Ԯ�s�(��kǿA�;/ŶUj��X�(�����X3���R�Sغ���u��KESϯ�%'���#b���0¦!�>g�3s�M�6���tŧ[��'QXaH=NVj)�
}���A��a7z���N���m��aH%u��# ��l��z�4�z�Sr(}���3��2�g�H}Bs�w�L�W��nθ:|t�:	p	��5]�˟���nW�V��L]E�E�u��(?vAW�J�ǿ���[���P(ͅIVޟ����^({��}f�(g�rg��5��Y�+��;Yd7��s�bu'_zAa�d��7n�.�n������^쟟P�q�m	s�:�@|�,�K��ST���YJ➓I(��u�H��g��7�}�j�c�T	���F�(U�<��F^|`�~��))�"�����Y������!`�\�o�cwvnhx2��-r47{��S�/m���=]j�]���d�%M%)�f�q�O���	I�9�|䆢Md���	�G�M��q3K׋�����e�**�,i-з������f5L�B����ZqxϦۈ�|�'_<u��Z���tR}��}��4�f�ѧ:�Q����8IIJP���f�s����ԳE�N��۷o������ۧ��V;��P�� .��gUd�x`�+���g��\�Vy�x��jN��<o.�~�{`�5��v�'��)d�^Nn>�������8�ݺ��z��٠��~<�)�x�"x���~w��M�5�,tV'«��w)�Uq��-��qp������ �E�t�H��ڼ2�BV=Cѣ"%��L�k}��~���?��:Y~��Y�d!\R�@WƴB;"�㊵�(ʙ��GU�� �Ƌ�B-�7�("�^�q�ɹ/���O�Э��4��r[@�-�pl��RY�Y�X�l�Y���9�Tϥ��Fu�ڶ�ɫ�韺s��݇�+7Q6�*�4�Rh�D���'�nΫ@�.6�x3D`N���4ڪDo�v�5�_��f}��r��ڡ�F�͢���x<?&��T��i�����w��n	bE��pߊ�(�Љ�0��a���)�9a�c�h^��Ч*EH�P;-p_�?�!G2q�K*��4g��&*���I����JT6�?�	�ure��ό2�^�s� ���$����u�x�m�1.1��M%��{�@�k�ɘ���vV��=��?̉��6:�-�"[����Q����C�5ܖ�7�S�"M�(�j��F"��V鞣�5Z���s�
c�*h�Q勿~a� ��{��$�(>.q��ӢC>p������5�����|\�U� ��/���w�J��`X$ 4W�be��L�H��O��9ݜ��k3��^{���L�_j���s����C�(�T��Qӷ0z(��~��U.��nZ\�y ��E�SN������\���x��9B�~��_��f� �V�KQ�js�B���`���2	#��M���
�c�Ë�C�"�1j�5�g��a��|��_Ȃ����h�S݌��/��9�n�V���!D1X1�j7������s���3��>�X��C)� ���=��>u�4�F�{��1e���0�.ɐx��n(�ڠ� |h�c��c�/�J�(=��͵��h>-[���e�L(�Q)�Γ�Sx�G��%�,
2l���tNF̡R�y��W�ֳX4N��}�I���F��p�c��1:	@���RW�*)J���^N�e�Eֻ����^��D��=(��Zf���ѕ96J�"P�|�B�� ���qz�I���[���^�_�B���,����%7B�a˶��*nL���0���#�1�J�o�O�C�yֹ��f.M�q�G3}���R0���4�n�� �[�n/oA<H*�S�1��8Jv㼡h��a\{��n��H���$�l �}l��&� �ۏ?���`��H&�D8��ŭ���}y��{��:��%֫�Z_
����X�6򕁔���*f12���r���uk\x����������Y:�L�x'�R!�~�
A�{Cu	�[eh��qlD�����G!�\��h��.W��C>v`�}���Z�����%���+��1��G�Tb�|RӃr$������B��ۊ癲�l�V��D� �y4R���ٜ+Y?�Y{�5]EX���=�|!�"���_m���N9-��ςTe}�z��'��߿�X�f��%�b�2Ж��1�.�ML��J�\�i3u�u�A�m(+8-<�AA�c6$��֧�����k�$i2�E�|	]%2圛�`=�}/�֕�;U�ϨLm��۲8����:hrJ��.my.���-^ƹ�pi�P�e3�ěOf(�؈r�oa[�_�˟}\-�#O�w��L%��:�D��m)�4�X�gl=@���MAK�0�i��a�������&��u�e���*sZ����O��iaY%^���֝&kg_��N4���*�7i[�;q�y�|�%8��O��S�c�x���C��c�|a\y
 oCJS�SM�����\-"�t�q�6��$�W���!�ˈ���ae��)-	-���c��Pkj��_�WɈ%,[������(:���4�%�2n���p'��,�`�yR�
S��͂U��\��Y�=��L$��Q�UMA9���%0�Ƒ�2�?�3<�IRi }�B	�V�ɴ6s�;;�I�n�,>����,���L�������"����3.�7�F9�䚒!k+	N�!��A��<��:�E�~Cnm?g??�����ٽ�=7�{�l����!0�m�K�
�)��T��S�� �r�B+Qc؀�49�3�"˪��8�am8L��_:�A ��LrH^�h��(`Hy�Z������6�@_s�����:��Ȱp2@�N���i*�\� hXiN.�{����|�v�?�XH���P풴�iǈ�4��+Τ��d6�0|���GH�87~ͨ�o��b�TiΦ�Į��y�m���S��=�8�K
ݶ�|�~\ń�t���(NS��h���;!�V�гdV���q�ڥ��-����������F�� �U��Z�vM�x���#L��w�|&<�����ԏ�,&�5����&}���)�p4~����ܵ/5�\/Mė���"N����U�$���c���7��k����c��j��ؠh�*��Q؀���l��9������ձl�l/R����U[��>��-���=kh7�/j�:X�Y|%6gá���;�5ˮ�;o��?��i�t�{S���D߻t@c�l���c��������Rx��<83M�]��g�v�C�y�//�=��>�4�ss��6�������o&�����ˬ��mgƊ����|
&M%�N��e,�]�*�c7.�ONً��u��@W�M�z�z�ca�����Cr �X�[-�T�
�������<l�M2~���^��*0�/l��D�F�2��$-���JG~��~�.f��Mit�U*�C�P�؍��m��� p PT+m"/]���g�P��\Ѣ8D,���ޟ�p�аY�sx�(dWC��p���YO�fH]2���rNv6�[^������%z.N�_`��Ƈ�..�����O!�;��ç���������1o=H�hL�߉Ag���y$���J[-�(Oƫ4U�1����̙�o(K�G���"�,k9�[IU�|�-�!�� 5[�ϓ6��vd:�C��Uvi�(�&�P���?�5{*��b�r����GW +(������ra&�P�Y�H��?I[]�>zJ�l���D�@O�p5�����	���/��iNh����Mb���HS>�*��
�W�����^!_)�O�˗�l૖���Lr�{��|�{1L�|?�8���dXY�v�p�	�qH�[��F�{T��sJ��~u�x�ċ�p�<�{Dɏ�ȅ�l���'��ԚN�=˵�@r����4��R1�,�K:u�����q��qB��(����y���;��TXhv6����7�.��XV�d;* �P�ыm�|����o�m��U_��#:�5�`�O������W���-�چ$�M�kp�(����>��8��N3�z ��i����a�K�#��$x����I<I�k �?���.'�s��%�`�B�*��n������[G�u6�����E���2j]���-ͷ�����d] �۹��z鏅��C��-��J��?�]H T檲
צҥX��M��r���M��{w�\�����D�9���S��U�<����=�8����6yQD�����TG0���ڃZ��1���3Q�c�n:��!Q�v�#��b���QI��W�_Oy���-���0�nJ�բ��zj�%Q��@���_�`�2���A��&B�& �������ښ!P����@��^���߉����G�����F��E��I����&��n��IӔb�b�]�a4$��z����I,�Fgs�2�R-��a��.�⤨�އM:
�o�Q��5�.���������D2R�L0��zY�g ���Zf�޴�@@�0��5��k��TT5ϻ}����8W����
�"MꞦ q&×Z��]�3x����[K%д�w�m���U2�?�Nn��_�M���p�e�r\ԕ�Wi�#�q�g���w�������3$8ru
�u�8�d�_�z�/K�+Q�M���)|��݇5�f�;�7�b$�VE
��!8��JvsD9�Pb@���B��u$9PΘ_��Nə��lQB�l@� _�o���RΦ�s��-��Mҝf�C�{�,������ʎV,��3�%�x���F�/��8�Nvϑ�F��
��N��S]�l(��<��p�֓J;��F�������C��*�=A�T)�Z�����p�g<t��]���4i�&�IP�|5�?�dE{����T�3�Y�ޤ����Đ-x��O��o�������@�֧�	+��q�����17Q�85n�!���"{A�;�:u�5���t���(���ΐ�/@�P�T?�x`��y�Dp��+{>� �a�L��ք̴��ε8"������|e��1�AZg��4>`r@b%��'*��Gݮr�Dj�\���e�����<_�깵'�i�$�������fs�&f[�P�䚔��E�Yc�1�^�]��95�,�u�T����#2 H�z���B�*�ի�$,��{`�q������*�rɽWrވꄞr"o�����?K���$�?V;V���2��u������*�Nj�m��:�d�S'eC��j�Z�X���0,�{K�#��p3K�vйv�C{��9yJG�P����_��h��纩�.���Si&�'w��g��Ts�MX o�'�t��W\%t�v�y�lL ����.��n����]r�?xT%B�̹�.t��Z�]�=Q�e���'>I�+5��յK�k[;N[� w�W�ƈ�e�x������P��7Gv��6����I�+	�A桌I�=����y�%�	c�1���I�˵h"%a�Lw?��8݀��S�+D�
�P0e�w��:����` �?pH�K�f��C�oH�����r!���[�� $q��\��l��;De�G��6x�b.�V��b�
F���pOZH���cru��$�RՇ��Q���4�0h
�	:np��t��d�H 4nxBI���/�	����ÿ�;;�Xg���t[ ��Þ,�7a�W������5:���@^�&Q���!�-�z�ro74?��4��cY�$����b[!����||�:����q#��)��]��vզ5o���>ۆ���9���]�l�������A�6�G�P;�}>�\d)���yz�	&`az�MOy ��~EWfb_H ��5��k��M%̭l㙸��� ��ðL)]�ad�Km{�#v��/��pP؇��dD�7�+�.�f�.�A���sX��u~���K�.�C����~IT>w�ۋ
��Q�Y"G���p�;fc+���Q_���N�Np���XC�O'�"�r���>�w�i�y$g7Ϙ�����6��	�G��A�K0�GH��#�w�����}������M�v]kn�>s�x?��&�}�-��:�`Mʅ��Ƹ�n�I�P�&1`��k���8�,�IJQ@�ձ&ږG�� �����O�7h���𽂷A��QK�+�ȩ�\��~�\�&�!3j�v��i�M��~|zY;�E�P�\(`�m���d<�9F@�ց�[�|"{*Ѧl�[[�:�YH4��z�r__ڕ�.]��a����@L��]�CZD�M�g�N��v���v^ML*�x(��Hv��=��Y�``�ߩ�����uE�W��D������4��JX��;�v�=A�U�0\CL�Q���d�?J�d���!	␝⪴Ƅ��C�[�#�����A�ѫ�Dރ��t�t��E���g�@�f��^v��P׳y�6�!Qn�f H��;�vgjj@nS��Z�?��&������Se#�Q���Ԕ	�<X���sb^�r�+���&v/|~曆�L�aY���Q8�2$M%b�]�N������A��ɠ���k�^��gi)�'���3�&�C���jw+�L�$�z+i�P#�Niճ����D<K����q���J��D�wP��i[�E��.�������">g��s:H5��m�~��wl�*�R���(�s�c���Sf���jK�eK�U����Q�l+n��xϺQ��zU��Ԭ㏡o9\���\*f*�WL[*��L������I}�s(E�I���e|���ؕЁ���J�)���?�@F���mJ"�*��q�T=),�\e�W9��5y+� x��I,�w��.�6�ۅ��c�m��,��O����B��3�b�Պ��_���LJx
P��!@	9�{�K�ɛ��5��a�X�>W_�?܇NQ3�u��oc̋�P��@ڠ��|&MI�bTF�f^�h�L�3 /c�[��ܚ�<E��mi�]�ᕛlE�!s��!z=������������܆�J�10t^Y@>���@�Ƞ/{�(Cd�ݡz�tܗ,�{o��<�m�J��i���p��cq�l���TPe�ݭ �v��r��M�-�0�v)�ꆷ`y]z�D2vg�����B�S����D��J�/��n��rGX���������0�V��WyH��^B��d�Sl Φa�Z9�^(L�yC��w���!,�a��2h����~o�����W�\dk����)D����e�tIq�<�7�#:@Z�6�"xcF5#q�-��}8����lm�h� �z!��L�f�맰�j�1�r��d)�,��[ڱ������]�;�C�JM�r����3�j`�b֌��,޲�>�Y�a��B��rw��p��������S�@,�g�(%E��=h�ôuG��޻i��O��ѿ�⠪z��Z,���|`�uy	3�2��Y�I�W�JU������c�I'0
}$��KD��by{r�¼��\�����/��#��+��)��M�I�J6W^C��	%瀉NgKUD�K�]�bh�Og���"3���Yx/��3�D����;.T{�_G�"D���g��kOz����8�.l��f�ub�m��_O|q�M�j����Ϡ��Є5tfHߨF�O�jI�(׉�Wk�2÷ey�^�2kNW50��J� ,^����d	gw�uD���� ]n`"ϒ³�H�����~�;(kQ�Y�2��(X�irD
�ըC����̇����=P��Kj�`�C
��w�&)/���þ��kssC娈�#;�
���G�qz�\ϑ۰��[�[y�L��@u��v��<�1�rn}/��d�0��E�3b��
3� ި���r�q+	BBKܬ��'aH<�J2�9x�o�$�^��s�	t��`��O��hfjV��#[�0��B��¤}K��*�[�R�	��:f����`�/#9S���Zh�Ť�J�O$r��s�r��ݡQ�+l�iE��K$Qu(�	PU&��Zԛ�/���c%���^���$�X:L���?�ZJ���' N:��W�nB�M��P��2%�a:E*��@
�{�װ�v;Ph�)' *D�x�R�l��exY�
4�h�O�+r�����y�,�!��,L��Wc�Nr��k'��B�)�8���d�uA�q��O?{/�ۺ09<5��s��a.��`Z�9E� 8P����e�R��p��dl��� �el��8Ï��<�kQ�U/��w1btϜ0�%��� I�P�Ő�nC�Qhd�;�Uw���Ւ6��Oȴ�i�M��C�/U(n]V�d��ԑG���SH��ņd������d���~K���s�y���_�t61��~�7��[j��5�p#������"Lbb���+��w��:S�X`d��a$OSb�W���A/<���k����3}Т����u�nxbw?��d%���L. �����'�t*@�ϋ�Ԫ�:`������@p2��*T"�]��"��Ox>
X��˳%��&L�Mmj�~�������c7�!�Y�w�w���ۂ��E��N����'�g{��"�����y�ȸ�Y_DB��������R�;��f
r`(�|S�����س��#�����Dr�%��E+��J+�,;O ��i�k_��F.� �e�%���,&�$�(��m��W�%�STa�b���l&��+5���oǢ�`����A39�7�кN�L�HCې��<���#�#�,��;����>�Ȱ>���DAL�)cȪ3���< �?��'���K+����c˻�GNxK�w��#r�S�z��p�yn{��s�V�K`>�@��ֽixe�fm�� ���%�VE�$�oS�c���ut��Z�L͆�H�L�K�eѤ�&����ծ�d��]�2��@V��T��D��}��]�jy�+��#;en@�L���͉�%c�U�L�L���
��+D���ĥ�';È����.��
�;1t>�:M%���11����$���yD�ݓ1��r�4�λ;dt,���k��tc?�=�jI����v�Y�u�"�U*��,hq�M�֠�f���O����ij A�S�8�΁�6��V����д�t�{�����f2�}����ct�Ο� F|�)�.J��
&_�� �K1{���$B�5 �
�qT#8p��`<�4#�C�Ӵ�ͨ��v+a�Q�00�"�*�4y �+99|+2�Jp��SmL�$�ޘַ 
H�tL��Ip{����	�����pl`���n.��,A��z@�*���Q�Τ����������~x�K8ɱ
��d��8J%�t?Ic��FŽ��˔_(�9@U��U��G[���<ɦ����I��D&�b��
;��D\~��:�+�A8�^���@�������< �㚑:3��d7�@���M����ꫛ�/:�<b=_!`%�N0���a��S�l����}���A0�4�\~��$��=Ҷc�1��kv�S�v�t��+!o��a����/�c5�*�#����V�2�k,' ~�{��>��~�R��XNl�9��2��-���!���:� �JT�eW��7Z�ֺAwz	V�l�E�8�#܄Z������/	,d���,���ap��wU~~G{K��#�:1q2`���?�$� �����@�bCs8&'�@�@��lY��t~v����0d�s��!�,�_B�-A�N&0���P�uj����yX(����ZοrLW #E�Ԅ%ݏ���kF��pοjbN�U�}��0��WBh�񶺙ae���f�%ȫL���D.L?}h�1'ᬙm\�^�I��V`sBy�l�5��L�\�՝8p@�4��QV�pm���("~���Cw@@"�v��QA�׸[���NM���Ch�L޻EZ��:>�����ly߲e*�K��a��g4�8|�$��_�U�����c��-p�葒=×���!�Xc1V`s�3���9��40�;2����x�uy��4���`t�|��b	�� v#,�S������a���\~5���1fJ��Ӊ)[�g�e7��T�o���]�� r�`����s��N�z}h�'���������׿�JK��m�`���P	������
i^�>s-g)Ἢ�q*
��h3آK5YO7�VX�X�l)h��5t&��:�r�ɐ��«v�RxD[{�p�m`��Mb�ު�V�+3��d� ~�vhk�+:7|�B�B��	R4Vza;׌X���g��#��$Lm��TzBژ�.I��#����C�M��|B�l�ε��������E` ��c��b\��Vi{��4���d��^�d�^���"�MM���KO�K~�iz���	��@����{r^G�	��
����Z|T���p��k�| ��yϯ���d��%����c%��}^�R��*�jr�"���>�҉��5�Ó�u��>���I����QU�}��R��Ŝ[�C?.���dpa��~���[�Z��y�[����s������*r2>�x�1q}ʭw�C烈�v���_K����r��� F�`K�s�z���ڮ॰���&+���Ktȣ��6�@/�fY�L)eh��@�~�ߗ9���RX �̕#�h����E�f� ��NGv���� ~�a>��	����r�V����"�0�P��}=1c��D|�Ƙ�d�H������!��f�/�:܀�|�lHPltU8$[��V��+�������_g���6-��T`���uM<�X��{�~5�f8?�)@YSo�'�������h(�}^aˍ�yGV�A}Èə���N)��-c���6w�'��4$G���f��jVτ#e��%Y��mcH�DOL�+~����,��Uġ��;0���;p(km
��tM ����n�h+A�<�����}�N�����Ͳg»&KG���]T]b�>W��KZQ�s�ƼxzK��9*�^.�����J��d�q|������c$9� �;j��)M�Z����'G�dS����8?�?�ޅ���㧨B"�L�Y��*"�$�L0�Z����C�04��<���L����$����m�M~8��! +����<R�P�hl?{�x���*�H��|�6���p�RgT���>bB����3-w�������(�R[3n�u���c�~��E�R�ۯE�D�hh�Pᛷ��� ;���A����Q�_�0�OTH"o��k��	G���2~�Ÿk���2s\P	����	��'��{(N�̶F=�&�"yk�u��}��@|�e���H�*W����~V��e���$�e)������a��hD��:5|>���&�b���j�0���b��{[3�ǅ!���m+ϕ�ꡉ�T��"���^xXxD1rb!Yc�1o�w�����ɲ3�|{p�R=���r���ߴ��X|��HU�Jk��o��<H0yhf�H;&���gܝ���C�0'�yj��V�A�S�x���vR��X�i���9�*s���c3��ܱ���(�x��$�1u^�ͳ�)w!���i`��T��g��̀���j=�f��� �����9�4�,iL4���ɥ<y~%w����t�s�˸"�4x�7Q%V�yV�s��}a�AP_�B�U�y�#��]{=���+��Pܶ��1�1��9�`T̽�$��?��/���r�f�G	[Y����˶Gh�#��h��4��8��x���2��F���Y*�2^b�4��T\4G����8kl�tJ��\������F���\���׌��8�#Q��I�p��@_�܁�}�LbL��(�b}��$�Qrj�6�ލ�C��DU� �Z��3~@��/�N�z����o��at�J��|�,�=�$V�p-��<�&J��E��/Z�i-.g��b{wt�5��xs6t��w��4��k�^:	�8殈�IZi��U=Q�)%���%�T( �� k*Hw�O�8w��y�b߃л�U��E_�Y�F��,�˺9)^��g��C��)&r���0�n���eJ�bL�YKQm�p	��6�?gҚ���IJ��3`GA�q�&��	0u��@�#�Z�Hf���τE5�_u��Ns]m�	�o�Z�=�4%�Hm.Υ#ͤ#r@	ǜR�J?]�/W�u��t;L�e�/����~�� ������{��9�|׾нp�J��a5��]��T�;�s�號�ݱJ�w*�p(驉͟$�R	[�љg{��!�]�����np�Kg��'��g�].&8c�p�����Y���1gVѼ���L]Ѭ�OW�x�r�>�8i y��ɝ!Zx��jo�,�S��%�l�c[`ܭ+g�`��(�z�l~<�����1=�e�\|%:����c=��q ��~-z-K8��8�Z�Dw�֏�C�4��xP��D/���׷+\�� P�$j�����zkz?�|Y�b+T�geh�Iy�b�n�ċ��m���ٔ�����?F��R�S�#�A:��S�$�~�� �RK�W�\*��©.G�_�31Y�R?K�\�gʿp�*��6)̶�"ܥ�N�I�CK�*D�N� �.3��0�!5o�RWM�5��<d��	En��4ə�����d\^�}�^b��)���+�W"�N�ՙ�V���BZ9��Z�et�[�>uJ}��O�*�*z'N7ħې<}48%�9_�LўW����=�'�[��H'W� ����Ӫ��Vυ:�1�x3���.�R2�:~o�_�v���Qt�%͕���V�⢱�u2a�8o�'u�蘘l����mx�eNI�I1Z��d���6Ӭ�i�[w����8�I�/�?x��\8��z>:��qy��WI0������%��Ȱ��i��e���T�I�f<�`L_���S(`����A��y�Kɟ55=j�>��]a�j_��Kx�
�rLj�D�(�.R���Rjq@�9�Z�����|iLd2��3�V`���c7��fa9q��Yp�]0h��D��앬-��T���7į�
� ��/���+�[� {�a������j�~��t���ӱ-��㟈�uV���kt�L}���/�g��w �b�:/�<��+�n*,�	8t�pΈpy��߼�^O�U�KZ�T^.D�YO�����O�">�͏]�{��H�9�����c����P$�����&()x�F�+���˩��!���Jټ�
L��QP�@�L�N�~�5 ���z�Y{M��{�ӍH���"]DӁ����\�+��$� 4z6���qx�h}�N�����^��`��@|���hA��V1a�M��q���%�ߡM>Yaw����6P��O�͜��}-@���g���5\������J���P���V\��3K4z����V�'ȱ��r����d��9�s��tO���F��WB!Ңb,�v�b<���wN-�(,�FoϏh�ł����詝��'M� �c&��Yh�)��[\ =�o;��1����i�_N���p(�OK��Y0��e��2�?�c7�<��-��1����6̉|��ъ��0R��������7��#�d��ݴ�!Ę�61K�;_��Be�;�~<#4`��d�O�FѶ&u�e@&��D����ԫ�
0|�^r�V���%�~�����u~�_!��*�]T�.\|�c,F�KVM:�g���
�Dc�X�&o��[���u�=x�?%�z����q��Z�L������oL���m���}6Ua�K�����B�O�Ƅ�_������a��<E�]����#���u\_\i�݋�+-+���+�!��v�����F�9�����E����� �e+8�U��<���@�*DXե�T�.������ށ�4EY�o�qi	���;gfg�����G`n�����.�.�6�mu�^oɰ�8��%1��>?X�5��x'����O5��/C�P�N�3Aw�L.2GV.����
���^jmV
 �
v䂆���T�y�,��8�T_�nu|����6�d"�
_h��ZG���ܕL�L�>��n�>M��"�)�\�!z�HZa��1���4!�"�6���k�})������btP��M�z�vs���KP�uh���Pۓ�ݜ�Ck}m	�������,EdQ𧻓� ��{ߓR�&�\^ߠ&C>�_uT�}\�d�S�5tҭū��%f�!�'<e�����\��p�"���\���ľ&c<9�/4L�.g�(
�"i����RK�	n��@�U�� P/�7y�N,�ʫ��?C��⇵��!�-h߾@f8zXLrYg#�좐����tي�s�N���,�M��b��&��=c����Gٺ���?�Q���0傽��e��	+7 �,�LA���Y%2L�[���@��z(�`c�S̞*rz��Y���C8dv��
�u�HbE�����8.���0r��?�e�	7�O8K�`ݽŇ� Z��v�h�z��C7 �d�A����A3X1L	bPfʛ�����
�S�+?�K9w�����"EY�U?#�
"��eb�hǥ�c	Y����w��1S����b�3H��Р�-,k��G�4)�'�%̧�? !��95L�ݱ*��ajc��Zzh{]����l*2�y\E��x9#\�Τ�p���c�����:��1�y�h�g��D������I,��<z(�f�@�g�ˬ�[|BX��،'ė�T�3.>/<��h5𞻇Ui�}<d˨@�cH�Pu���םB��I�'pbF3s���>~Z\갡 �k��)��J�?��������IP\7ΘGX۵�.j�%�&pG�8\�B�{�I*��G����S�c��짭S_v��b'��A8���p�6x�}~����)��Uq�u룧���r#+�F��`A�ZlR����~&.�[ {�Zo0������ST�[������/r<��W�}�f0�:4��5�bRZ�օ�l�c@�v��Cdn���h�ꑑ
�<zM�9���h�P�:���e4z�r˓m .�g�Ϊ^� �t�غۦAQ�Up �4]n���4�}Gt��1UX��=2�>K��M��������c��z�r�?Fs;?�L^f"������s����ْ��5+�=(t�#)�Y6�`ME¢txG�R��U�݁PU!޾ܞ��g:?N_r]C/u%��)y���-�$���fj��s�Hj�<﯎O�G���I�j�@����*?~P֢�R�;�N�Q��I g<�:o���5ȫ���/�##uA�,N e�`6���{�L��P�'Y��,����.N�UCs�B>S���`'(��-9.ͥ��L,��1�O��:$����FY4�-���)\�o�8��o�0eE�r����X�%ɒ�벃�U��]-���G%�u�>/����[@x����(ՈB���(ҹ�=M�l�;�k\d�T�o[1���ɸ<�>X��ځz���J��`بOw�j줧//�������H�0�S龉
H�4a�M'ۛ�fIg��s`���[ٔs�\Wu�r�hdZV����j�Tr��ssR���j�z���O�9�HL���&�K��M�"�Px����e�7[[S��[WD��[���X38�t˄�s��戡.�f��(�_&��b���~O+�e������cɆL?��s
�؁;��5;S�Ș�F`�}����(�I=\�s) �<S����Ğ��Cޫf,p�o��֠�H��޽'{]���^, {IU�g>$n�nZ牢 \�ʟ��lc�D��ܮ,�Y ����z�_A�`>���Y(��7^��f�?�� e;$܆��Q�e�����P���&u?{*��6{#�*�L����{�Y��JAH�w��}��<W��_�^��'g�TZ���}Y�#F ��
�e���* ��LS7��T��mJxT��JA���K�<�/�6��&i���ܚeU����]�9��Hَ�z�6i����?�5{|�p�?�.@u���)�S�1`dB^,�_r|9O\��5�'���.y
�cg�Xv�@�?Qg#�ё�*�8Ry�*��A�(�];�HJe�w�د �~�C4c��rIpi�ot�k\�?���>�'C� j��c��z��6DK�+DdƏsZ��mT�]k�X8��*t���Ԃn�V��C�~�9��g�]�#LA ���{c�|ņ/�J�tu��N5��C8�n�n�!O��q[cn��Q��1���D�=׫�5��S����^�@su�$s�p�55�|�
E�C �a��3�3����/�_ZO�6�5XJ��G���>[��; �NkHj�t����Xkܚ�ʝ��Kc㏲Umm��v�a����:V]rh���.�"I?�pn���`�+�T�֙�1�⩄ݧ�@��;��X��5#gNW��*���n�l�� F6"
J�g��������Z��
^���M0�r��+��$���W�Q___J̠ic�\R�<���m��q�K���"�zU���S4}��Q��&㏟��!��ڿ} �6�
����:r )i��{�U�ZS����O<f&_n{�Jc��#�гk�ۙ&�<�GϝI����~TU���Z��
��=b^ۋD�z딼�YhQu�:���s{�!"F�� M"w�3�b��3j���5�!D�[�&�@��wT��� �ߋ�M1
;7�Fվy���l�������]�:��2��,J5�+53� y��s�	��\��$�|
�yb����Q�f�������u4Y忲P�ƾ�x��8��l�<��`�,���t�c�L�$ߥ�_�<��,9���}r��>3�y.���a7�d��l	yXŌ�N&V��W�yv%�0��EF���`k�e���ݎ��#�g\$|�4�ʄ�n�_9$@��:ckxe��د=|ą㑐�#����K�r�c��戶��W b�kD�/�,�W|�����>�Yh7�"�UɔLH!@Ǉ���w*c�*ϧ-X����v���a��0��fke@��zb��oH�!�a"� d�En��Q{�~(�i2��u�$� �]��j��~��zǝw��ٳ�� �|���ڰ�����L���ƅe�R�"�TW�H�62Yo��2�v_���)�a�i��';�9�Ƚ2vL1��N϶H���.�p}�)�1}�Q�����m�[������/O�&�G�(���_�'9��:�ߕ�\�+�]�Z2����դ�)5��0z\l�	6��6v�6�_#E߷(�%MM�1��vN�T�)����#G��Y��>Ǔ�f�+�\Ѽ�+�s����st���Hޥx��7K �����2���g�e����;B�,�L�}�����$3{x���$��Zy�i����J���feu�x!@{�x�4�ҵ�;0��ˢ'�������g��H͔��>���@�0����S��N�O�z���œ�?��L~��¥f�>a^�`�y�r����RE�Z��X^!������CͣS��Y[���*�������	8?'J9���b�}sĜ&� uB�Læd�U���䖿�ϖc沞��;�20��������`��������X�7�Dy���Q���Nz>��~�{��R�3�-�Dl�挤�����4/v�����,��,
�'��F��9Jm�e��^U̮���J<���a>�i�Չ3SA�9p�]���s.��1�pU��"5.�c+���O@��\/昲�s��*��R�8^�%DYG���$C��ү��0�uт�����QD��i�e��	�i�dW��rrz|-;��'y�D%@l��	��8R@A������I�#��oF�k�N���7��� ��n
�}R߱S����M���ˉM>$�'��7F-��M���Y�����"U��&�>��䝰�潔|S�4�%�6�;W� �0��:��q�S�}�9sb$�h�8=l|��qHCf�z��0U�KGN ���]|o����h6��!��S�[��ryڶ0�̾�LJ�ٌ�4����=��VҸ��h���f=�F�`����1����93z�U��A�x�L�l�8_3^*���fi��;v�ة�Ok��{r��@��W�G1�)c�v�+�c�#�xx�{��6����:����JfA����%�����s�Z��( "��I��������m��8)����r�p՜����8"(��Ö��ⶫ?{�]i�q�PT����ĳ��7)J,������,Pn��X�/�A+�X���qux�~���Ӑ��ae�թp��﷕�L�Kv���sU�bG:�㷇�"�+��}�+�X�fM����
�)Ķ�m�PQ��U��Q��}F*=���oe�i��}����>�WVF,��*���2_�/8�pU�|���O�|I4!"WB�X� N]��IB�Ȓw��Pk�L�>��8K:'�wjś��=�dp{V.x��/���-�ó��&2���_C�}�
���b�ըV�P�F&q'g�h�%����2D1e)>�������)�BIIc ������5?C.���3��S��P�i���4ss�y��;4ȉ���Ԕ���?���I���N��WCqCq!Ȓ�:��A���`&�N<�(�	S0hѰ ��bM�t,J�Q' �=cҷ�>ќ�^�poF~�����~���|�-�gnP=�����3�]e����O�xA��q7&&u]��>&7��+�Ҥ.��U�g7w�4S�.Q_����F+8���g��G4\�^�x�Idw��&�y��Òm�Ü�W���r�i��ӧ0�G⼣m�)�}�B�X���gO�����4VV�Ώj�X�7��n>6Y��o����}��#	6����<���MI������)�L�U\#O3�'أ��!ϲޤt)^E}�O�
֐��Ĭ�iG����i?�yz�;e��z7�6�{��q���[Il8���%R�\tiy�G�fzg�'�p:��3Vl8�<q����"��ɤ6�mԅ�R��mN^��Ss�f��2��Ogߝ�%�Iם���a@�8q��#&�h_8�͒s>��942.�J����S��2]b`�ۉ����H�8Ug����u�f�@��Ի�au��"p��F��ep�K2�鮓�Ϩ~��d�-x�$��4�˦��ba^y��>�`a�_�H��ס	)��U�xw��nٰ:�3:�N���=��!�
د�z�¦|�b�.ZE��nlW
M_V(Z�s:)o-��VF��{��GP�����7�r�����1�;kc� ��e��ܢ�/��P6:s�o�g,D�=�"I�">�o�F�]<�E���U�)0<Z>DO�X�FN�U�nYo=Q��E3;��� ꨼��A���"�;&� dX)��<KBN-M���i�����cI���P�\o�]#�#����{峮��X��s&��E�zv�.�ZQ`-�ո��c	]jH[
ls��1ܧ���0�(�.\�(]s�X	�.�v��t�m����n��Z��|��Jo���i�%"�!��49X{!��c�?�pm3�\�;���$��<�1�|�w��~�jk������⹘�\�i)2ɥO-�IK�	�RZ�Z?�%�~X�ԅB����it>��e+W�rk�	��I�(푿�7��ټ<Se�LH2��(���h.>�tT\��;\�g ����*d�Ŏ�׸���`kVB!�Qco�0W�i�>]9X#`����=e-�\f �0�^#����h<؀0���(nd��<)/T�f:�L�����	F	h`�o�կ��W��B){����厪?�O�������'[��< �%��\�q�+�!2/e�L\��m�അ�O��94��{�!�L�{𞬿��3�B����-m�uW�R��g�}��U��N��ٵKQ*⒁�p߃�2��t������ @0��[Z��o����W�����k��1��b�>_�w����<耵��6��S_�NaL(:ch�̎���3�G�pF�1Z��'xbǝ�;�}���"���Z�;S�-��ɍ�,��� �M� �����z�eI"Ѧ�|�
�sF��ع�A*�Xm:����c�T��ş��̊#�)���J�w�L�_���L�
�;��Ʊ2J��&:;e�52o$IT�,�Q}ޯ�#`O��� �t��j�E�\���m4AX�"/n�J��ik�i�Q�R?�:�bt�0�Ɍ�^��=��Ж�E��8�Ռ�����lH��� 6
��YKF�!jD)��pHa-!���~=K�I7�$��`�5�p�Td��Ԃ�0�M1�X;d`�*ν8u����iIMh�X�����r�=e�ܬ�}=#�/��K���7�Z�	�Hn{L5n�eA����ThZ?]����O@�V��J]4�;��z�9���(�(�n��b<�>f(���p�P�X�lV�藴���O�Ǳ���Q�u	.��A�2j&JAǯd!��<�IyQ���vͰ�ʮ��⍵n���������4�ӑ��M�8��4^N������X�݆i���������T�"RENS��$+(�hwB�O!)~������Z���w�d��/�Bk��]�l�b�A�0AOUo��Y�̦�����+��Q$!��B\�>�iB.�i��f�K#y�9�0/��bjPy�n�|$9k�S�}M���ق�_d�
�_�v�%نE=���K�3�'�����#� �RI�H�7귖�.��3���-��D#�/��!{�ڎ�QR�7���?1%�g��s��Q�=_c�]�L�jȢ"RM�L$��>����ʑ���qf���/ɺ�g��ux�R� ~l�����(��:���!��ger#�; _�a��q�֙+�Ѓ�?֜�u۞3O6I\EZ�"@�+W 	�~ju� ۲v`.o%_h���o�;U��@<�D�T�����g䏅Ȼ
�c����,"��u*<�C��P�I�M�6Ġl5�g}G�>����!�G�`8��ظ��!>P�q���1j�<�8�V�9�Zxz�� c|�oC��g/PutŸaƄ���j6�1Q�t�TU`/;g$��=����籄����?����
�Tm��к'�O�f�1��S5SA@�R!f�����;=1F	s����!�2_4bm̤��'�F͛,�h��l�y���iO�+k�Ĕ�!�A,!�Հ���O}<R,m�`xt�8s���Sa�	Th�FDu���7�����m�����!�H^����v�9b�eY�]f�����
���9AW��Y�����7Ҟ>�h��K.h����.��ސu ���q~ ���q�
�0
?��!G�<o�����pz�T�:�_'7��XO�7߬� Sl.�/<��d�x`����W_��� �{aH�So+�ʦ7V���=�O�UG!�DC��;�2�̰�b�ó[U�KEY�>�)2s��ol�J���Y�:ͅi\�؂�X�����6�D%Y�3_���^��<��n/�Δ�-�Ԓ�ޛ���]��e� �R<F;1�i�ΈNx"AЫ��d���t�X���'ק��C�d�Q�j5/�ĲBs.�m#M���_��]�y�N�O	j(�y*rH�9�t/D>/������`���/	h�D>:z����er*����_�$A@�{�	`-)�Ź���Fwyc��:�)ȉ��!p�mY<��Wi1�X���z�dx�_5K,E�i࢘���DTx\L�D'�eQ���v�d����H�jaHoK�`'}Jd��!�U��32��p����"ﺌ�5����s�ÙA��ˮH�����*��!�#����v�~�>��Z��6���w3��	��I4"��#UH�"��d�;��vw�В&���ʭ���.��(y\a�P4���E;}f<$�������UnAJaS���[(��6�M��"��|�w[��,�L���g-��`�@A�F �t�b�;^�IK�˱�y7a��nߊ�:�M��3��b�a[�[tW O#r-�L�G5E��Y7miͣ�s.A��9&��tY���g�L���
�DQJf�1��z���a�r�	��~YN���[m�U"�GR�mf-�3��mՃ��؛���##����k��yU{��'R��.�� ����&8=�{c��$P��~L"�!��m��B$����Z��;)���Ѵ���抇5_Q<z�9�a��(���$�tԒ�{E*��2�s�pi�"��K���iLB�	J>�ȓa�����?"�W��x揲'�����1V��az�G��!}!��褉��],�[-Ni������ S\V�Sl���Q��C{��!���6 ��9�ID��I�&� -p���f�ň��c}�dQ�-=�V|XA����@����JLbT��K�f�<p�%��Q���s뺣���T+?w_���P��`�H��jԐ:C�Sc���٥#�tRZ�g���p.���K�3!kmAw$ۍ&�mF���e8�;"vg��ؾ�G�%/-�*w�r{�\��Sm�Z����LVA�p��7]6F�QҪ�� jX����.13���]X�l�@�����D-��& 0et�I����92=R*���)�����뒞9�o	�'�M�E��|Γ�K�ă��9�Ee��ƌ1`����C;+���M�
��{�T^��e����rJ*��F�2}l��zG�����JմGWqo����k�:�q�;�}.�A�(�\�
��,Eq�?Y:U��A6��y{������^���E�>�w�d�
�Dױ�0-),�����U�00�#[� ��������8;���yl��E�o����x��Q����Cqu !��i��mT1U����-C��xR����S������E�C�ɂ��Y)ဴ�5�H��iX�&#�·V�G�x3y��y%�\��|�#����Ð���2�B2ȕ@�WS�A�;���Yu������T`G{$����K�ȫJ:��;����N�ȡ�κ�c9�����$�a8���1�*7X\g�gq.�9�村2'�G����M����"M\��r�����MJ���р&r�ԕ�M{ܗ�W�`��Q6Fm?G6O��p�i���"��.�YD��F�z��]�.�	��e�;NT���i�,�+���w)�|2��)�_��/��Rvcxd�&V	�V���gҎ��^�.��Z�M�L�5ǡ�<��.�rj��X��ʻ��D2�j��eA��:���ݬ�_�p/���V8���Z��Q� ���%�_��ҿ�6����[Ό��Q���i�ۓr�n��<UT�RGyƣw�x)�H"PA�X(��<i)�9-n��De�	U �͈�6M��'Ap�M9M�sLg��b˘��te�,=V����Ɍ��,�NRbu�H��B^��֓M'�_B�/'�7���v��no0���%�d�� �W7"��$M��X��9|"^�{S�^�4��]o4B��/3��:	�1��d��`1͐"�7 �5[J�[�jW���I��W��`�EdVRS�ie�"?��t���KǲMl��4�^��i�'Q�Wn0$�6;�W�%��R�� ��}Y;�4[������)6.zꕬ�������^1���/�
�^)� cW�����)U񪿘
N�&4�4��>w�k�FQ���,���aì%�g�JV)"\�C���������'rؗ�["l�7-�f�j�,W�a`��잕��J�g.:��έ�dD/�.���
�#����F�L\�X��9����蔂�G)���B	J��jZ ���\�q�}�-�0g��/{�
���1B��lI{����_�5l��d0�\�����1��L�d�+ƴ���D�]�D�};<
qZ[]�����cevӨ"��M�	Ѭ$󧫲ilC�C�����,�%�!do�\�@0�b'/u�ov����1
|:�*�GU�4.V BmP�g�g�0��x�XE�s�ٙ���ɚ���������.��z�oi�?�_��K<αq�8,;�r�&H�7��V�4�lĩq^���a�hO�K��SH����M�%s���H#4����d���[�s�٬A2�4WE�>�qrr��Y�2�C�Ff�����-
�|�m��h,7[�� i�:�ސ��J�[����+E�ύ=�P->��l� 'd�,�{�{�x���Q�Y�gbN��V���g�����p�Sc�>�I�����4��zk�`��������{=7#ϕ&�r�j)xn�8<��|W�7�~�3���U��-�ŘO�e�=;�r��p�ce8�
��G��m��;�;26�QM:�z�� tq=��R�Yk7צ�(X��Ɇ�����v���<�����	έ�SX!�e�=�9�Y,3����y��g�7�"֒�Fy�ɗ�4i�MK*�'C����Q�DiT�{��;w�J��z�s���պ*owp^�'{J��
�g�k���d�oI����];��C����n�1�vܜ�>��܀9a�G�]�TW�F��-�{�4��%>�ʫ���J���v������2��+l0$�!`���3I'8RJ�|?��/��2#Q��U��3��.A}���Y�t��٢��QlWv�����WAO�(�o{��O�/�^�B0�wc�ĦA�XV�1kH?��ag�J��4���;w=��f[L��pr�PzyD%���f�+�s�\�F!�/�K�w<�Ou�"f�{�r8x��!�V(�Y���?���.t�P_ U�'C�a`�T��}{^=#�&�?��?��������r�M��%:b(` c+$�E��z傄`0=2�e��4��;ŵ�P\�.�ߥ �@<� �v��TD��J���&�@#p�ex.}E1"h�E�}��y ����A��Gbq���_?=/�e�LJ�՟T0ov�4�S�ƙF����C�J̚�nް�FO��6�=�ZEȚ0Y�R�4��!ȫ>y��ҕ��[�O�d��޺�����Q�dn�i(�Tut=Ռhk����j�n��hd�(_aM���-���ܚ^���=�X��?@�:Bq�%�t��0��U�a�ڕ8[.�� �m_rpL������I?��1W�m�`k���^���/�����b����dkS�����U<B�*��TiF�����<���_j�}a�ET�E��Jw��]m�^N�݂o�����{�F�u���=��9[EYd���ռ|v�@��s��� R��X��b���\�7>�\�֜��@[�#���;K�<�~���+�r�x�����.d=���⺩�M�j6�w�]6"�HF��|�T��ө2ňX�5hR!�T�5}�TEh>e�I�m*���Yd�vY�Q8zBZ)0����Z7�7yy�&�R��I�<�����E5�-���^+�gQD󗶰}P�=����Ӯ�Ԡ��_V2� B9���H[��qN���s�Ŧ�r䧩�vb*������ɲ5[c z��_�0��5��*�qUVu����QcD��e=5�5�����P)�(�ɱ�=�,�-:���$�O���8�j��i��aꭢ�])�J.U�9��
�?@��&�v�����D&͡x̓�%g!$��ո�i��-5���;P;�1&E'����!ܔ��Z�\��\>R]��F���6U�����.ה�S^B�N���I?WQ�9�ж��s�ؾ?�z�l^�[Is�n	�798�3���h����&��A���ɐGYP�#� ���XNϿ�!�_[�=�}��%O q-��k�������^ң(Ty9�3�`�kX�f;eFa�i�'�mȍ�SL�9�ϋ�N��7�I��k��p����|{T���m�@��������bKlkACiH�w���F����͏��S�"4b��#��̤$�a[�YYE��:���<5�=S:�?G ^�������=��dY_x:��4l��.)�Y����ǗH۽0�J�n���.˵M7j,���,
hJ9[��Hu(�QuU���FħX�a���#�<��rz��[ �'i�Be�W�a� W&68iG�V���fL#�Z����
�����Cz\ϛ
h���-*sE�Yp6AKh���9��5�#�i0��£2¿UO%�����qi��b�1,vZ�xi�nΘ)8�0C�":��TG�J� g����sq�xو©?���
���a�+��y'Tu�)�.���>Q5'����"��G�����_�{��[��=�z2�h�]��}����ekh.�?�E�D�GS�5�FYΐ&��{r��ֺPx�@]r��dˢ�_b;�o'���ϡ9t�������X����zR6���򖢸��e�P�41w�pc5�6��ng�
) �@�T2ߥ,En�ug	�\!��(N�%��r��a�t�I���Mҧ�kn &{|��;1�[T=��l�M����ݻd!�Y�M��+6Z��Γ�-������3I�_Qv�7�W�[�5��������Ar`�z9���d)83(�Q�����q}�}��i�xg�P_�ȫ�#�.k�_i��6��>��������_�Zb"��M���AţJ$Xqf$����d�9��ײ�F������9i4g�	���� 
ʝz���y_�p�i��a��<L��6��	T��o$P���	=�-�V��n�t7��|D�2(n�kt0u/n{7��E?0n�$? ��9�R���9Xݑn�g��o�OaҐ��m�k����LE�f�"�D���RN��1�����__��A=<�"*�Sݭ���U�����i���~�y�֧�g�pzp��b�8i��%6mQϚ�/a�%_�k�d}�	T����.�ګ�4��[�I�zC���q�J��o���@|��o�?(�U��[[�F����u�i�	��W{SX;w���cY#�*�VWY�֥tpz�����_Q���I�b�����.��	���`��ڲ�8!�u�QK�E�Q����wԟ�����]��7J�-�֕!�+ŕg��`v*�"G9����Q?̼f��c!C��I����Y6�8�9�v��`���G��K��5K'R�bY���E�I��/0}�d[�2�ҡ��2 ��cr{^�/���g���
�6e�}?�PW}8 �%lC	@������cϋÅ��g���W���@�L%��@����"��S�0��[���}�H���љ�C4��?3܃W��ؕ��qt���n�e(ǽ��(J·�f2	 �I��_Z?.+ gy�3�ˑ�~�dk�hM�$��+E���J��KC\�{(�k��b�a�ӟ �%���c$�X���}��D@wsP0"�T�(�P&S(��@���0�4
c� �4C-Wω`譺w���q���K�.�Ls���}>aA�I��� �h�@h"�"�n<��.��H�����=�9�����be�,�UйpNCO�b�{��h�p��,���j���|�� "�bR>^������]j9"Q�Lo�����nq�����>c�4?�~�S�F�y�aU� �"��������[�.M��j�kD�������հW����k�l<��6��Jp9�츥��V�Y����9��A|���v��mRe�m}4�$^1�
!��O�>�a����l��)e�U�����s���̩�s���@Ke��	�L+%�#�R�Q�G�����[���;jwFP��/����S��E�]�����P}����}>%���#�P���hd�7t{��)ZO>t���O��f/
�
�'͍&�L���Qr9��Y;���A�⊌k��������nI�0�L\� 0��Q��R����HGߖsK�/!��~H˱4@W4����� �l/����>xq��0|���N�,��1~b���W�ξ����{�G�
p�lX�&�1�YR{}�S�h��l�
",�ӡ-�8�Oȁ&R&a�5rV���h������2����h��lI��F/qf��w��-p�G}�����ۀb|����	�i��;�f�����Fh�){|"E��,a��![��y ������Бr���q
[B�\AE��8f���C�� b��K���J^x�B�
��\�5��5W�c$F�F��p�,�P������[62��d!j�l�]	����"��
�r�`��Q^ �4���xeն����������tӟ@�1O��v
B�c�A�!�����%�m��#��>amA��Y*�a�ݵ:�4�nG��{��\�2�a�x�G���n��t��&��mFr��!�,�x���k7�+#K̃7��"Q8�<D�3T�����X՚_I�8 �U�-����;.I}���ɋ�F��-쳗��������&�S�xϊr��?��%�^������w�Ȗ�[B�]�@��X�*�Q@��F��/�6������D5֩h�����-���y��%{���{%��Ћ}����I�t@��	'04�FjyRe^c��5_���[�v�C��t�J�Z`yu����3u��A�(O%�S�AA�G>A�2����`W")�n���P�ܯHP���kЍ�ʴۊ���],k�I��g%��g�i@�h�wƏ���l�2n����DL����� ������W�&^P,��S���7v�;X���w�n%�aܙt�ߗ��� �ݕ�yҊ��R�0'j��9��T~~�������n��4R���N���ٞ����i���"�eF�����݉�o��-��I$s}�����GF{�qX��/��y��D\o�ρ�$ڱC*@݊,{�hǆ c[�]@U�hUTXߵOF�ܣt���0�[����R��D�̈ 6�+�|Km�di��sT�>�s$���1�M��.O��S�_�p&���k�e����.��Ϟ����Ɣmϖ%�nF�*�>|g��2��q�Cv� Mg�h\�V~͉�T
���������"]�j >���I�cc�UgV�uӰ����u�赍��a��79A��3�l��ϲ��,y����]�I�m|�t�F�@�pή�W��-}��q�xqr7�8��z�x���#�D�K� ?Y�Xó�h,]D�}H�m��K˖�|)�>֡s����~�h2a�|��_��<�Ɲ�о�`|.UJ�+�:�� �I��&ڴg�!uf�;�ʮ�0��a��3SONk��`
��T�*${4Mޑ��Q#C6�h�Ԋ�e�"�Ϝ�N���>��L�D�N��-	C�� �w�5	��
Z<���:xIP�� �CF�yʎR�KT�	.����V�MK�
�n'̴� 0�����/8O��Kڃ�t��#�~����m����Ŧa
��c>XG�uG��\ԗ��3(��W>�\R�U���D(�Sn��ej��%�T>� ��b��Y&�S���� �9Oﭨ���!/}����"CV������(��e'��jY�&��Z'��a�"�.k�co�N��-��|vQ��@���fL�
n�$]��P�0�"j]��V���!�Y_��7҆���j�J]�\����]Ӫ6��y�t���2%�'/���EC�� �,�Z�jǣ\@*��"�?�o �y���M�Z��&8t���0��1H�L�
�^7�!&kPL	�c�Fr��~Ә��!�|����^I��[�Bh���|%�h�y�F�򛘡�T oB`��xKBN^�Ld�ׇPP�%�7P�W���R����*S>/l"���S���y�9ZB��O!���y���qZ+��hq��pK��N�����,�e��2A��a*N���{�$*���R�����9R��Xߓ�Z�� $P21{��ĩ���U!���Z�s`�8� 9� C!6abn��5���'�Y��Uw�Q(:0����=�����	)G�`��[Y\��2Z#3��&�pH͚
e�hڞ��y���W*Ϲ��<^��t'���PS�wO������H�~���E�i�4�D]j�ϪA���3�:u�ss�O�PѺ����~�\�o�ߒ�s�1���
"
PR�V1Լ�7c�(A���hK/p�O��)��g
236{OM�S��#Z=�ckcY��qC�6��^_QZ@��!FwU�tKUo��Jj�v�i��|�_�#�K�6�~�#��,�[�\H�!hc?pm����`���g&]�ti��v9ĸ=¥
)�k����l0!��5�8%�5�|�+���)@����]�t�A��{2j�Y� ���|������Z��2�J�U�8��Y�G"��Hofu'�t�Ff�
�C�|H�kKr3��i-9��� U&�8T��������^̆	j��A���N-�����}�<V@l��*`$��y����/�FE���!�;�����O�NE�{�'��n1�M��A *��m�~>n|@�*�>�g7�2���d]�ȫ}/ʛT����̑�g�N(kKO����X��1T�9�����l��F�������2N�U�V�%st,<pȅ������b��*e�0#�KPo�l�c��Q�H�K�M�������}q4Se�J]gl0q@vS���!y1{��PMݡ��>�2�7�<'e�ѽ�t�Aߍ�)��Qs���>�>�:}̚'
%�:�Ѫ���{#���8"%�&���a�S:�\/�F����o������zjz���!��r�g�7>w��䏙3$��7���Om��|a��O���
�w=p�������x/��LH��x�����1I�� r�=�=���}�\�L�HgBs@�^��uhm�ÀC��4��)&��>���ǟc1�Ӑ�����,�Jn+��I�Y�W�΃�I�9�
�% A��yr�e}���w��S��H#�v����\8:�F�U~v����b�����u�(�H��w�g�M�]��pട�|Y*4�sCU�`���2+.0e2��?�\hJ��aA��.��t�]#��6�����a��AT?���bр���!
P{q��i�k��A���^�����x�}���g��j������t�.%#��P�I�Y(�*`1����pu('6飙f��kk�Ѽl%u^���&�'mԞ�>O��F@�	$�l�4�+�:����);p����������x�n�mG��=���k���!0�|�O�Es���-��SU�&$��i�.����ӈ��R��$Z�B����qL=��T�I������6���"p��EuDr'_�io�j�ٚr������0��w4A�1�!H�����qᴴ�b���A���ŅGc��>e$�S�pqn���A�m���o\�eDuf�^ �tX��]y��c�v�ˀpC*���	'��\v�2(o�Vy ��&󝦮U��`�B��{M5vV�%�ʢ[@���D��U�a�욤a;��L�l�7A8�8�t���2o�/�f޺p*����=`�.��x�#��<�<����9s�+%��(���7n(a�ϊq�߭������׊�M��y�g*��y�I��~
�L���g]�O*A��b�c-�*8W'��P������frϙ����B=KD$-��-m_�������b�c������Μ��1u��r���G��ƺ�{�T١$t���*�&��7����������1����S_}=������7<֓W����p�B���G�;d��b	]�0=�4��c�m�A2Xqv����Ə9��)h�FF�?��9Hg����ٸ,�/�����Lʤ�:sW�!���OE����+�d�jA���,�N!�,~57��i/ʠ��;MMǋ�凲Cl�ɶ�˅Bl�����-2(o_Iǳ�tQq}�O:Î!�.X�c�Є|EYu�duG4��:�M��J��Y��E�n�/��RiC�ܻ(�)y�������[�U��Z]�Y`������T�C���f����b����F5>+"f���.�����U���'|Qh��V6�%`8�Y /?L¼,�#�O4�ۺM��9(��M.��K�Lbe�bp�� 9fey��^[%�������@r���8/�+�r�ц���{��5N��!g�܇a����3vb[�3(w�~��;��=��1Oqd.I��_ꕢT��]i�q�am�G����vw�ޔ>�8R�J���8=���1�(&�JѠOݑ�P�Z��ٱ���.�V�L�,��(��j��/հ=�c:^J奙�0��v'e��}4�0+-B�%�ҙ���d���& ��\�[M�^PO��|!P��U�:dɡM�d��P�)�7l>oE���L9��F��簟X> A��&7ݬ�s�gm����_��X>���ƺ�O5��s��(�V�������ý�?�Fp9���h��_��?�P��Ҹ�{>\Y�%��#��+2EqRc-���2�h>
b*�����\/<5�׶�lʗ �W�_:�⑷Of�n͏$����?p���%Yx7�'ړ�EqudA�+�xR��?���Xssx hރ�����S��k��3�����41!ײ�bd��6Xܟ��*1��z��O��7´
��*��T��̧z�ɒV�ۃ"�c�8�ߛ�R�<����<g��\��s�M����=[�H4�ќ�y~Q�a�x������q9m+/�3P����>��O�7��O��N4Q�V�IVkG~��֠�n@�d���TB���$A�p�,s,�"������j|�k�I%�?�/L�+#�R	�x�I�-R]@J�䪣ܵXa-���;LyƇ��x3���$^;I��\�� &;�"�1o���d�W��Χ�ڇ����R���}I_��E�)Ţb�>��haG���|���c��k���j|5����i�y9F:��,ͨ�F��G�&���GRn�j$��C~�C�u����C�)��9�� �l�����M���R� $&&��!�t�|M�] ������*J��Z��a�l������X�|t���s�ψ��|~�����Tt*�����Fϥc��N��ߵ���	"�W!�jd+�b;!Uz���j�A�sn���Ҹ����h�-�h5��/{3ھiAh��w�g�`Fq�+]u#�;�ƅR��_pz�yM)ȡ�O���A�d}�;�2/j"�v4�}3����M��;=zx��qP��H���E�3�<�(x�yZ }}$K���|}������[�]͔~�t�ƱCEM��I)�G�PJ�=�n)T�40c���Bߺ 4��Q��D��P�'�O]Y��\fs YfkKR\�Ks�0�X�V�b�H���I�zi;0�-i:��y� h��ƌC��$u�������v����KV��F�Ǌ����w�z5J�\��m�Q��I��ԡ߅�c�}H5�Çn��;1{�u���O}��j�Y&�#a�q`�{��t{��/��|�Y�� ه�Ƕ6=���$@�be�{����af����	���W���Ɵ�Ǝ�Q�'�bK�q�&ap�l{��9ZcO4on!Z�W(�*�����۸+҇T�m*���F#.�k �♥�}����[�R��U�x���<�u2�͔�T5�d�2��G��,0�s��q�S��d�F]lHՔ�~�����u�C�}G�xv,vp��_�: 	.�CH���H�-�c�.���T3^��ޕu���{濃��Nu.�Lߗ�ذ�&0Kד������N�E�i�YX>��%c��7�(�:�CW.�>E�5�=K�����6��e�e ��ݵ"�UH�p��U�����;Q�x�ٚ�-ѿVh�w��caG�P;H9W%rêP}��u���C�e���k�O#��<�<���/t��!+O4v�~c֟l0x>���z���Uܪ��c��pH��E�wNj�#��̋ܚW�!2���Y����Hl�`C�59��B`u�jhCB]8�����l^��:�
�&�CM�����	��{���� ޱf� ��!q���%
��Ms�������'OzO|��>;u�{�h�u�	C!$����Ɛ��Ý)Mu2@�����!�c*MUs���W�5u�>�,I�k���<C�x&z��#�����?� ���
nI��d�f�� ���l�
f�ԇ=�>m�l^�ihC��IDfň�����Y!1O]��	X��9`$\еE�4����������/��=��A��A����&�o�Ro����~���Gxqsq�V�B��f�p2�:��!�������&|���U�.�hْ�(�rb6ey�ii`#8��yΛ7�rr�9��2�(#����@?g9P`�����e�IO���X�3C!��q�ii�πW܉X�v�t$��4�o�,m���7��ku X�����>�x�7Q���L}6����B�T�<�7$�����Ƅhu �&?�	E=�����g)0�R��P=R1H3~���-_`w�v�cS%Z�_��N����+�jy �N�3lƈ6h{�� w=�� -b��H+�M�\�eöN瀙8��Č� $ �p��Ч�Ο�]������O]K<Svm����sbB;Iur�`q�Yz��%S�̤���k8 fM���0\N*=�D����2����Ж����h�ի��Ry��t8Q������ kK�����=	J�g�S�q�h`Fz��4õ�_NV�ӿ#+�8h�_��� c�S�N�>��H�y0��}�>�ꗀA�����I��Z���?k�Cw9��6����r�F���V��1S���D&�I���:L9i`�i�D%���}�z��->}�Ȳȡ���:l#1_�+:ΒoH�pwD�b�x�@��>�x��@�/e�����u�f��!�C�&v�ӊ�jU&З������l}��C_��,��m�ѷ��Io��H-X6ኺ#��Y��{]
�z+�p���@�ɻ�j��?��4D���� R�z����n6(�)��#,ix뮊+����<��`�D�⛼�hH�����Ѱ����ݬ� �?k�	��Yaq�«|=��7����9V���l�mQX���x�B�9������?!�D�	�l�[�w� �AI��׋,�J�x�=&Av�b<�]WƘ� �Ҹ��̈�O+��ߧ�
���Y÷����0�b[<:3�+uj�ls�-,��򄔭t��ɺU�Q�9v��7�f���B���[Z�	e�2�6
�PC"���)��5��!�}b9�J�t�]�؎\Bk�iI*���җ�dųܨ3.�������qw�]^�FyKm-�Zp�$fpǙ�K�L��_{~�&�vj�G�ӫG�N���fօ�ű]$����U�9��#H>�r��`�Lԝ!#�Џ�f���4���?@P�X�{�{j�/�I ����e}eH���U �}B
 �R2�!���9C��L����p����I����������y��)�]�H�|�#��A#��u������XG�cn��sx�e��ma�e�5�~�@^F�Zf���J3i�r�����	�:a�v�+(��JL�v���7�،# ����fr$NCi��G���݊���B+(jnh�ew`_��mЋH.G�
�<C�������T���}�q�6͋G��Q`s0�\��;�0�VՅ�����Ɇ�IV�X������g�I��U;�^7J*�q:bO{�\�����K\h�Y�+��B�"��Y���p�\�}RХG]㒨;N("P"2Ӆ����F%�h	m�D��`�)_��4���Q1���A�KѽR�?�ƥ�s��_y��ށJ��p!k�Կ�U[_C1T�Gc��Yл�}�����G��� ��nZh9��
0������}��.oo\~h�o�")�*l.?T1j3U�|���W�FӯMrj��c��w��gaθ�mev���c�o6��:�B�@?���˲��l�}2�h�<}�8������3�Nmt��N�TɠCD��R����k&1Ս�zA��=
Շ��!pC�ʂPq
����Y����i�[�.���ʙ��.��������7��jk�؅���$k��"d�pj�"]m���%r뗸���������V�B��g��z���l�����
$5�nI|!Q��,�����a�D�92^\	�Kퟷ����g6sUT�vs�W�PtiT����~���f!��ۃ��9�v�|?�s�!Ą�{���xe����7����y��?-��z�Q�~R3>�����qmQ\����T��]��ĦyՌm�j��t]z{�h��E@R���D�s���*PMXO;vk#����g0�E�@��֧�̄�Oe@�*W^�]�}Y��Ft��#8*M=�q�����t��ݳ�4is`Ԇ��ӓ��� }�k�����(uD���V�ҩf$��\\�j��bN�@�d���.{�c����X�Rjݗ�j(@��-%h�4�)eg!.C)/ó&qzO�"cˁأ��k����^�k����@�-��׵�d���m�=��V�m+&+���ɕ��jֆ6����Sk͚���=V�Cv��[Ȩ��̛[n��p�ΌK�u �i�!�K�(U$u�|�51q� !��~̚C*B��1�c�i�n�E�-�-�վ�JGX��1��.f[�T�ɔ���˿?��������~,�~@�09/��|�q'l�:r�JQ�C��O� .g4�g���<��Q�6'�6~����ڜE숛Q��QYLDh�	�����Cw����(��ؖM� Z��������:���7���|�jm}-�5�}�]��&X����{�s:����@;���/Ă9��m�qh?�c�I_��~��pu^��&Pd�wma����WՖ~Ʋm�t*D�ȻP�I��G>��*�
���B��V��oX�@{7�Kh���/�ڹ�Q��w 9WZ�	�Ev�7���f�X��%�̊7���:��#PC�2��!OM��p�k�zƊ�_�j�v+���ne���S�0}w�����j���ļ�q/8;+,b|�Lza�*xUS�-
��v��)�DrD�$� +�G� ��E2O �)+�n��6H$�lby�-ͧ�"H� K]�F#m�Wv\�8�A��]B+��d�۔ ɓWtQ?I/���g4/pj:hEVf���ՙZ���<`�9��5�؁��xn!dk�h�hԹ�_ޒc����d(f6�M|ӝ뀫�e:���PaL�J6��8o��b-kK��8=)�l_�N����<�!� NVa����y��ϐ��FEt���N��(�ZQ���ZN&��ze��/�1�I���N��)��ȏ�7vqw��'�p6�%Q��3���5-�����Խ��:	h�V�.F�0��d�V��6��-l� '�.�Vy��A� v���H���`qo�"+��-���D��s��&/?A�g�x���QE�}z�$�olKg\��>��	����t��=�/u�A��J�=��Kj�#@��y�4���d�g�n���v��'N�Ȑ}�cv,��/�[ip����QxMp�2@�-�S �6
��B���d�,*C�6�i�w�vEp{��g��C	]�*�6�M��.g����v�B:�x��^���U.�Kr��}$L]n��.�7$+���8x�����3�ub��Ӫ�8ʀ�K�t�`�7�hWM�^��K�)�#C��(=a$�F,p��+�XiKj���H_�胩;ʐ�@��n�rU5�f�[�����&��}g|q��oI$�s!,uAa��t���g�ήs��HD�\�V�]��t ���q���?��Zt%x����XK0��q�{�ş��{���
�
=�^5Љ�q(d/�
Q�H�����Q8��Z���'��e)���Q݄�Ӹ$�"z�q��&
09��,eu�2�}:'ij�nW�������<Z�,|�b�x-u�ܠ-_��9���&� [�F���(0�J]�1�@�|r�ÝRS��,~�/�F�F�����v����q�l:��!�:�0k�a��������݉�P����LRf]�{�鼳yo#��E�xd)�(�;�_��<vH~T�1��O�\E._7r}'�}D/�D�1H�|]��a�`q����	�9�Q �i�b�����������q1:-���:�^����&������i�|�.|�&Zx5h�G4$D�m�_0���+���/'f0a}r��G��y����z��<mgɇ�A���7slf{B�RnP,4U�	X»��Ú�rIY7�'�"2=UnL�_م����4 ������P���%m$�����pB5u�y�?���4�����{���0A����=��w?ф�R�^��d(ʭz��k9����L�D?�Z����Wg�kx
�����9�3�뻂���YMK�E���d�R��\}x>|<�6���>I����kF ��Ծu��� ��h���\I��`�ŵ�uQ
Wd�G:'֫��R[�l��@
N;����G��n��f�B�P�O�<V���D���a�����g����x퓈��{g |��Ȫ'����|%tm�h�C��rE����[�������Ty��4��F���u9���I���A��5^%���3 )f�t�$�Ha�ƀ����r_=��1�x&�v���^ÈF�S@�yo�)@�؏21���u��i���\ϓY�|�?�v���^�t30݌�Z=�F����d�OJ\f�;M�^h�lw�f��Jaz{�:���S��Q���z�)�{���<�<A[,$�C�IC�{^�Q7m���>Wҹ@��0ɽ��s�\�w�b|�5�>iŁss�9pE%��ي�����5|[���
�O܁�Tw�.��ڕ�M�#���u�4KJ�	�����y���'�8�9���o"�W-`t�3�"$3I����J�h4�m�x6<�aU�l�t��Y
��)Y������kx�4Z> t�c�c�(��?�x ;YF��G6�"㰵�>^hP���0��{�~������W�׆f>Ӫ䃾�#$�~m��Z)(>��0M,��|f:!�ϳ8� �������7�ϒr���*4��=y���D�Q�'���ȏ+
޳�r�r����z�D�hX~X�� �	��R���+
�w��1R�]9���ĘoY~�Y1$9Iy�51���Zo��g��xjC$4��ʠ�L��1IE��J��W w�e��� ʕJ⏬�4������?����x�Wwo�z\��.M��?E�4}Y�t-���2������~��� ^JԎX0��3��LKo�+� �5񹧼}��R����;�Վ��>����p�0[d4�`�QA�Xp>�e-����0<�#����(�sq�H_Ų4$�Ϻ<҂�%���!��fXs��&��URЕ�{��� ���d�����*.��Dv�NB�R�VV��i$[�/y��n̖�,f��a,���1~��x�1�#��di���_�7���r�ܤ��ݲ�Y��hR*Ķy��Ʉ�)��g|�+�t���)���������U�G���21����;5�`�s��5��Y�qu*$�6��?2�3��Q��N��Jf�/[��l#��Vo���1�uq�E<}��)��q�˯��g�Ʋ���{��zM�7�ae���@M�)K9w�LL����)d�0?�= �5IL�W����whY����#��`n�:2G��i�.��rq������7d�V ���Xwu�vF�qj�9��Wo;�������n� YG/�|����s'��JM�f��P��رc����.*U�@�Y,q]��v�7�N="�����Vڐw�!�N]<��֭o���.I�-���_���9�,�^�����̝���H�;��jX�Z��7�*Zs�Z��Vn���4iΩ�4!W�yE��h�����USR��=s�WS*
�u[)L��,��p������{�:���d���Rr1���%�
-I�l%�F��@�m�0/�l�a��H�+�yjR���
�D��D7�0Rw������p��,-"�"�����2�!r$��=�d���u�r�)�e�a厰lC��?�c�d/��\[�=B��t{�i�ܻ�4�GJ���I�z$���T;�'������C�E�}=f��n+~�H��Q��2�\�w+he�e|��bo�x�2���/�p���Si����tټ�$a��du3^q�x�F�9���:`GMd�X,,9�ә������ZKݴ,�Qǡ]Ҋ;���F6������ԩ�[U!$��UL)#���m!¼���� �����iC�/�b��ԪFn�Ү�:��aߤ"f����~5��聻, Lu��,�v�P[���
5��42����j-�����%�1�{F)]�p�gx�H�HJ��V�_N?s�߽U�����e��[�����_"��ۚ��fkX�f��n����D���Wf/Y���E=M�;���P@�m]j�2<-�s2bce�	�1������$~i�?�u6i�b���׷�0�$��{�nv��e}kv��2����Ƞ'�4F�q/��9\��/2QVA��,��t�棸M���S�A�f}�f�
 e��b�n.���/�ދ1i`!jIL�/�+����i4���K���j���C�׃�9Z-�|c���^UN�F&�Fv��ßW�Y�M�p��_<A�BH��)�~(�h[3�]Y��*��P�;[�qT�%����l�F��������n���0�^63���V�e��I������ˮ��&I�\�}�v7�ù��E��v5;��|]܃����w<�z�i ����]�Z���"�2����pTFn��!)@#�?)��a$��j�l��o����]C�= ��5�EZ|�kݼ*�` ���&4��eY�h�}y��_�M�+lܼ�Wg�����!Ta��K�w��+Ri�l�V�W;���D�Ou�s�������~��S>��a�z�Dw���+��D�䡤��#�ֹ�nv�ov��%vc���h:�����Ҟ��=��8u��D�ARkP69ռ�$�6��5)��s��qD����X4���#
�SK4/����	ug`�|��̕!OsC�@��S���������`��|0#��ܸ7��4���j�f������A��2�GX�����~�>�,*�$d�F��ϯؤ��f.oQ�\�`@A�G�ٴ$J47!��Ը�A5��׽;��-��dF�t�]9t��;6T쇞����R9�ƌp�P�<b������t�y�����$�� � o
�쭭��2(ncd^?��"u��I!��2��6ghzO@Tx4�۴z��e�wV����?L冉��=���/��M̋Ȃl!�KL�.:G&AƧ��:�-�������O���e:��\H� eQyx��L�_b�rb���݆�E�nX}���kƧC�
}7��6����o���i�m3�"Д���KO��Ԉh�$c���I��ɘ��egٵ\��y{��I\�� �2���{���+\,����
�@2IE���zHo��D�=�|9���^K��"�y\���<T%t�> ��&�LX�9&�������#"���j�~��o�^�|��O�k7�f�L����f��-~�#��e�9��4���7��F�G��M?����:V�H
��j�6"h�pN��(�U���ˇ:_����3�w�/`s�sL�<|#<$������w,��Y&��`����-ak���pq�T0�@;u&<ϥ��~/|��#�&\���O���[�G���x�t4E7�D����W�^X/ԋP^ql�r�����x�\ J��ta�F�?
&��k���&��U?(o`�Z�/�[� Ź�Q�O��Ⱦ�嵎����V_�n��o{Ô׮��K�P$C���0D��?��m�wDb/�c'~��kӒ���M( <�O��Q�$�B×�a���,|t&���i�ZЂSR�TT���^�xg�-r��S�2n��́��HNA��6�~���b I�x��|��7��I��з�o�,"R���%B���u�޴��EYλ��n5̵��6�ֿD�J)�l|/x�/n[�f��3��w�O�+F|�_?p��vL�4��3��V��t+�t�y�5�������Q�ރS�{5�l��Q��ya��I���j���߫	���Lt���f�xXE�N��c7�J����z3��^&��\��ga���OQ);~!x���9��M���7��n�� � 0�dC��Cy9�09tN$��o}�d&�P�3�DU>��)q�,O�K�u���T�~�b�n�q�N�iP̮�%�R�%�"��H�6l5|?U{̂��w�{:x��0�2>�Ue���7�+M]d��N�T�	=X��jpI�X�h}�����ߌ���pp��jd�O�����ɍ,45B ޹S�ߩ��z7?O���%]�Cyzx�1�e��w�X��2K�W>�,���⍄���y�3}����:�(Ϋ}�ݎj.6�����.�;�H}�5x7o�!ȑk%�	��!^	�}���+����a8S�1��㗏�u�n�Y���/?J+[խ�x2��w�8��(�v=;�X�)gg�C�S_�e�P�V���v����FUV˛����u���=��/��� k�!�łs�jc�3����.��ſ����-
�/1!�,٪��� ������Bˠ�� y��an�F�O����/�b� y!-�e_!8�#s�+�	���DJ�-8SSɋ����K������'lm���H�(��KP!:旯h6B'����# c��HK�5Z��f��h�K��iې��`͗cD:�>��\�V����fD�3�k��4x�%5��~�S'�t�\��0]l�K^���+%� $��F��ӂ��������N��D����HF��Ѣ{i~:i��.z{����0��j�nF�u�U�|"O읇��=D�R�og7���w�R:-^6�Q�=j����Zk����,��)���v�3�9�~~�%��-���{�������Р0
��´Qvmg���bZ����<���z�E�2H`�]
(���v�q�oi�..�a󇞼YnӲ��[��:׎2�_Y�� �/L�0>h=��*9������/�������`��R����?Qص0�Y�j�VX�bR�����>�^� �����GC�Gk�˫7U��� ���1 G�S
�S��ѿ�ǣ&�gpr����\m�������6d�y�p|��_V��;������u�$��L�:�*������d82� ��k��cC�r�l��-�R�P����#Sr��C`��>����vq��}�,��_>6dG6	���y�ү������~]�����C֜�|8h�H� ��)܎"�:b!nt#�*�(�v������J�Sn��>3��v��?֯ڀT9�]@�c�w�g�mil�&d��T~���bQ�2/�f[���hyf������2�x�UQh�\�{�d��3I���[CCnSڥ���]+�� �%�W�y��&J��~Z���'12/�@x��3P1}�dW�w��9)Qc"��h���ښ}=�<ri�Ā=t �t(:�r�ʖ�v���oJ8��=��72���1��;w藔~ёn�勜��4�,�V�f\����$�	}��V�XSV���a��jP�L`ĕ�l �\s��/�jo@�� _��l�
�KD��Q�k�3�F�<��{Oa��/��&�r�쵥�xCe/�%�b/��T�.�37ǥ�!0 ���!����rq��̄�����b{6z�uu�5T�F�8���]���79cw^Дl���xx&��E�����g� sW[�$�"�d�I�G_�l��'��xuP���k-]5��ؑ��P�����"��0�b�t'�yU��������g�"�O�jv@��_Qޜ<6��%L�A�d��u��v,�7�F:K���?�d����
U��ob��.Dy�(]�'\	G�{�xX˦/�|��ig�o�d�-v0S�!Xqt��:SҼ�ڠ�-b%\?�40��Cy�kw���΅X~esYF�f�_�	֌K�K��*+7��ӷ�����^�X��F�����F+.v6�&�sk�e. E�����x�jʎ�^�>QDѱ߂>���v�N�Z�-'���51c����oo|�,��S|13�)�Ps�;;^LM8���蔉`�!֞�iĊ�5�a��f�[��q������Ćܐ�m�O��: U8淏��E�t���c_yJb����$���Ǌi��F�����KL<�`��.J�P��i�j���IT�|��K�Z�u�����A�c�i%�$�ݍv���oK���%H�^*�N.���$�"p3n���r�G����������e����*����k�g��P>�wd���Yt�dx��4c��-�6$�%¯������8\�L@�&�5B�� "���W��,�̈¡3h�b��@�p�����Is�~�ʑ�Aj_���tH�4��Jm��jCac��+sp�rf��*<{��Fa���;���h��C^R*�Z�dwPOF�B�goJ#x�
��ia�97^��V�\y���\��$Q�	a��l�E�U�)ß�&��D&P8��w�g�[=��]I��W�]�mQ�E� ��*����fZ�e��)�%=��󝼆�+F1� �hxƄ��f0~H���w��wHH�3��~ѷ�2�c���׋Nw�k��4�|��f���]�������䆍鬅O~Q�hxn]׀��F����+N���@��z�����OK�͐~ѐәm{2�-�Ji^�EZJ�J:o��#Qrb2�3�,G�K�~m3v���_O;��xP�Wm|�I��?(Qd�L�T���:���vz�uY���?�Ua�J,j̱���=������,$���#���ꍉD�O.d���R���&�O�n ��+�ƔZ^�h�f	��tV�\3�?U�C�=��ǮרI=���@]g�*tv�WG�)�
mL���ڧ�IP�a�z*���6�XrT�7`��[����q�nC�K�'��T|�b=z��E�����Zr���f�����_pZ�5� ����Ĥ?h�N*͡��B��B����$�	���-�͛H�Y`y(�� �3�4T�l���hN,�'!�v)^HL�(�;���5VT�YM��p�����1��a��UQA
��(:`5-�.�I"E�A�]<�͆��u�c�A�ys�{B�ɦ:}��L��*��_�QVl��π�w$�lU�~Xy%!�ꖁ	f�H%��)��,
)��ۗ�3`0U�x��3�J��L��9�G�a
�O'�v1�����>��I�:�Q��0z�)!��#��$tgheR���3ȡ 4O���+d&��R.jI��"	(��&�\�
EWJ\5���0K���%{�^����ļA��r��T�%�_�ɝ�ו!m.�@�T�H٭�.�.��BF�N1����`�1�i�I�ړP�|@R�m���rq4B��e�AC��"����-�
Gޭ�A��],vr
rǢ}� SW��.aW�<��D�vGD�V�<3E�Ҙ�s�X[t��[n�0�K��$��y�� ���Q�~7B��b;fL�T�_��z`S��T���ZW�׊S/�҇:r۵_��}+�ف	+��˂���j�3��^�������^�m��]D&.�(y%Bs�Q������@������z
�	�j�:W������qw� �m#/L�c�O��Es}՟�$���ʾ�*^��\����F�v�P�a����3�W+h%�m܊x�k.�p��zc��K;���,�tYӼ���'<׸�������Uܨ�T�s��F�&�b4�p.�0=UY� ��"�`�q�y'�u��Z��D�G�Y	�?��R}(�y4�h�͆6Y��R*�dt�"}��~/Ֆ�NR�H���>��Zq�� "����\�o�hAH{4~�-]�b���q���W�/!.�!�|O7���և%�eR��+q��Ra�Rρ ����fb�(*�.�a�5������F�khy{r,p�q�Y)4FQ���s����#h+]"h�N�2T��3g@�Q��z{�� �U	xG����w��Z�@��=V���\����,�t��k]aּQXb�?��M%��p�e}H�fﭝ��3�`$+���⛜�Ձ�j,��&�t;R%(���hk��i}WI1����j̿��d�Fy�� 횆����HJ�5�܍!C�ꠕsL�6����vC�b���0�;�D�;�T�v��0�1������q{tT��eO)p,��S�6���퇙N�Sm����Wh��h)�?ʽ�8Y3�7�� JJ���vX�������:Ls��0��C@Jכ��/��gی�"g��?U9�_*9��;s� ���}7ss"��g$��F|�d��߉O�	dVG1|o�m�:q�#���o�¹��7�
g� �I'3f��/X�������X��RG�@M5�&������]�N车j�O��P=)��k4�h
6a�4��g�3xbY��S�C��ہ�'M��Pby��$�I�[�=�jc<�7[埩!�/�l{��T�z��2p\\9�'Y��xJ�*3�������	[�QU�i��!/J˩pZ�1<�+sM42_U�a�i��	�X"I�����Ψy���e"$�M�,�����C����JR?�c�+@$�WU�,�� �H�g����i�׫	pC���0,5I��H�41\�vA,�a@�I0��9���&�q=�J~�?D�C�B�׹���>��ra�<h�f3�6g����;t��R#���>�Qʴ��7ݿ{�m�����2����D��f�ߤ/o�|QN#$0�h�������>h�̢!���:jì�g�\#?�I�|�}��Z������v�p�^b/����s���iS`�у~ݯ?��.^�):�O���r��J;&�M�������I,v�{��<ј���6�m�w3h[_d�ܽ&�m������ b̶�h���,��q��@$�U�N��V�w�`9�ғ�M�\!�2���1���
FƂg�P�w����T��H���3"�q�?���,��pE�fm��fo�M�s�v�#G�lT���^�E�� ��6V8�|}����U	������D@�꫶����/��8��ln���F�������t�H�h��'k�X�D�tT�T1�-[���������S}O��x��Ύ�3u�n�;!�-/;d��҃�@���T�q����n�\�=o�����a�2zCf��9���Τ|��z�̋
0�c�
����ȃx�)i7�O;�H( ��{�py0׵"Ts\���G�c�2��E��@q��{��5`�"����(3�/@����)P�C��ZN�?���(���,(����Q�	ה�%�C��=�nC���gR��T�r�+hmL]/��y
�<�"'�Q�g}mCB��lO��:!|���\�ְ��>���|������R�ά�1>��S�?[��z�YN�@ % /�' ���v��ސh��j��C�|+�#��ṩ�"���75)��*�	�g���I.��Y�+uBj�v�I�L)mH�E؁�s��?�k2G� "�`�)a�{���|�x��WPK��QHx�Ѧ��dv{����TgamY�5+����ŵn�9���4@���&iB��i����	g�C�2����\37N���%����R(�)Ѯ$����`���[���Jܢ��^�����G����aѼaxp8��pSt�2q
�e�0S6lT4}-c
�T��pȴ,P?�0S���k_��z(9�O��p�]�dX��ile��BZ���G~�<�	s(�R�o�ItpU54 FU�՘2h�U��
#��cE�&�d��{��o� I��'��#��W��s���Vx�U�~�ř�U�(�9�;(j��TU�InY}S��+ef�&��@�L�Tݹ��ޚ;Aq�Bٌ��Z���e��D���~ۅޗP�=���%E�`m� �@Cq���3p]^�/�Ha�O$g�Sݢ�'҂sf�6>��߈Nx�Χ����H�jvK�h�	�r�㜃/��^SE;c���i]E$��+����{�F��ɦ���?��#{�׻�䱅���A'v��.b���uc08~�������=|���WB�U���-4`�w�JD�є�G�2���ӑ��?�i�38�QX	�2�[��}|�#���H�.!�M�Ό/����n|��)��BK,� O�s\d4����Vsj���4�Ni ��07&����cЪ�L�q�z=��(`�"笩�R�.�	8݃��X�աR�`�W���dJdSL�z����� :�8���e6u=n�9��� ���M��^3�J�W���^C��Hf��@���A��w��
R�����)x�F��մVfa������Z~�ͫ��d|�8�������c�0u�&�De�������-Ka/�E��<�fj��Ws@�����#`��v��h��x/�hK�$�q��3hU���Q��E؝��.8q���zY�����<�5Z́�5��]bSr^>���1B�j�LL&6թ��p~!^�sT��'�;��~g-'g�5,l�"�k� xcm5�:;&�Z,��z�ӎ$�M�g�	�!/YQ�\#҃�|aV)ta�F�W&uy�rA��_�#��"L�6
��wU(J^����2�ֵ{�{��O���3G2��#����q.�~jxۼ���j
�������**#\f_��6�M��!�.�E�"Bz_[�ɸ_�����c��tR��1�{m7���x��Aazj�����eI��玨��A�qцJ}σ���%�{*�էJ�*�¥�m�3���<�4x���8��y�)o=��O�gx��lҙD2��wp��U����]�7ӷYY���b�rj�'�k��IkC��t���&�T�g(FJ��L秾3���a�@a��	� �R�ךv��4���O���X����v������Kpp ��]����D�-Vm2�f��v`^D�*��o��7۝�;�n,�1�mn6b�:f��e!�$�;E��Z^�U?Y�$03�R��bm��{n���j3��5���tu����@��#P�<��@�S�XFSm(y�h$�qt��;\�����ۭ�ˉ�q^'�J�(C�;�	����BE�4J��l�/<�4���U�4dw$,� �*T�t����I��{�F�������+L�u
�/3q�D� �����ꉕ,�7�^�ʺmD,w����{P;3?/�S�t %�6���ER�w ��c�p����x��,��+EY$�߁�HM��3w�����,c����36n�s���y(�<|!�k"�Lp��m^�:M�
eC�
�:��o �:�-�-�@D�-H�-&����V��m��C�:����X
2vUo�7�V4vX�!oi�����W$J��
nr���:��������Sތ+����-6��*.�(�l,/V��-�� #%fTr���S+fޔ�>�����S���/P�E%"�cZ.2��3j�B�i_��}�qFx���8��Zz�H�P0�!����GG���oUd"
�tw1J�:l����58Q5��ڮX���� U�����D�xRʸ��'F�8�bf���S.)����u h莺"K���TE-RQ�-����� J�>�-V�v���h#��I2�X���?����aN2����p��#���
;}���������8�mN� �D��+9'�[�\TQL���4�9��7�ϗ�Ʒ_��ۮ�ɑ�z �ay<��?b�Q��.�M���\���:������ �;�)�52Xy��/4'6m hQ�^m�� �q`k�Σ�pN��-"`�NP��փϝ-�Ŋt,�/���ޫT���3�\�1�2 �ܺ�0{黂��x�%�1���_���́.��K�I�P�HEvl��dv�1]�k�7}zWėC������&�{�d�l:q�U\���q��JYfXr���z��~�K�W	O��C�[{V���L2e��$n����d�Ԭ@4�3b|5���Y3�A�>Z����w�T�c͉�ϝ��W�8:d�g�Â�!��T�vA���6�@�s:�z�;�N=.���D�$XZ~2��f��LEP�?ʷ�h7:��
����'Ղ�p/g�}k��J��O&���4�䡀�{+��؉L�t�_Z�.89��)��n9|�\��z �Y66�d�p� �݄$J�z1yo��u�!��j]> <O�;+�����׉,e=g=������4v��.F�N�s�'yEh�� g@�ZS��QP8�>��oHI���E��@#���	�b��(�H��s0���L�'O-�^�s�tc����-ocp��H� �������aE�ʕ������b���I�������-�OwOJ���wt��ߤ��wD�(��}���H���R�Z�VO��`��:y���c��R�J0���mU���%F��v��a�R6R��)�s])ů@�:�|�eW�R8f<�����d*h��9p�e������������V��{��Ր����M�Gi��3��M����������q��W��tb�:S_/z��s\�J|E�=8�h�q�F�%jL�6j�VlV2���#g��۲�hp�9E��u-�Z�[1��x�գP_jKk�N�\�.���5B��p��-���q�E�|������+)RH�W���H�n/�!!Ŭ��6j~O��tB~�	h����TBMJAsh$�Ui�'+n#�zٷ��,י�[�$7l��U�� �'���!��ݞ�f��֠��Jhx@�&���b�܆��D�V��(�ǔ��0%�� �V���b��y��%��ʽ��t�z+&���h�KFk�Z�0�f���-<�Q0��p�k�|?Z�}0y�_2k`��Q�z�~�ιΣ���'Kc<�rkK%zS1����}"I�����:C�ۈ��9�����oz��#�P�Q�W8 y��S,�L��4*�D�#�g��n\Ve����/��u)��e��g�wu�xp ���|.�����IO��
'.6�W��XXQ���憫��)���c72M?�h��(~����N5��Y=���I��f9!@^����"�C�~�Ka�G��1v�~���G*�\p9�<x^o�=��p�v&:�o�p[z�l������Ī��"Lߧ���4�6�[<�z'\���"+B�����f�� 4p<6�,�u�!�W	}�Q��+��_�hxe�J1yǀ�f}
~�������N��}��J΀��%����:ˎ��˕P}�^��5��ȹ�S���y��i3{�b3I�`�^�n��v�{��+��Mt7\����T��Edȿ#׻H�$��z�s���[4j���{W;�)9:����[a��uJ�L�ok���| ָ��_D�bF�B�Q�U:l�នѽ�D d���O,�67�O�0�ޘG�|�TJ,u���4���x4M���Yð�Ʊ�9<�'+��w)ɿ�ូ+4Z�^�&A_%,2�����p@���}�	2�m�ٔ�J�m� ������ji��ܖ:�+"��2(}�<��DY����	d��>'"S8ү�>�)wj���<ѲL�x˻_�y�B�苢��Gm��hTӔ�q�8t��O����.^����%!O>��Ðv���h�m�$�%B��
R_�{���Q	9����B��6K+�;b�o����f�?�r��%��Y#�C�� ���.�.Ϝ��[Y������u
H �)$,L'#W�`-�T=+1@8�O�_y~)����p�@�_��;����j��8i;��T������sb���+!�V�]F<���l?NO;�r�g,$CKL_L�<;_]�X|}@ضF[�y��������ĳ���������N����7/�h��=�޴gbB��HP7����C������ƿȁ�V�2~`j�^o%6>v~��}ҫ��&y{`M���Gf�%��u42�]ǹm�d������V��֔�]�A߼;pe{��sv�׭KcyMP�0JLwz}Ә��};^n����<����y�z�#Y���$�*�+;���/9p�}�`� ���y	�/�&��h������d�<8�J;֡�Yr��wc�?5�guL�.S�!�����	���9oJ�?h�;�B����"��pT��S
<�(n2�n4����K��*��~��Qչ�R�k��`G���S�a�/6W9��T��S	�o���B����l���w�}6���uf�h�}�8"{0�?��a4h �7H$ʯ5`Qw%	s�����; u:���r��X���%2�����TOR�1��GQ�ύ4H��.@�N���W\E����}�'M�1���q�N2-�2��q��'�M���� � �
����5US8���<E��*�3�*n�������K����1d3��2O��H�6�

��~'��Bc�
|u�Y2e	��1f����:c93�%Dά�m�z)	�)őL��b nw��AO}�&@�N��ٛ��|�~ΖU%�"��GWJ�V��2���/z��*���(3��8��,�4�2��n��G���Т��;��N�dX���QZ��J&%����sc`5a������}u]�y ݰ������iUm�r�;�Z�u�]�ƞ�p�v?+�|W���Ё�m�8�C��bo��H�U�^;��_�$�m���j�l�J���ă?͑�C��b,y�#Hp���&�m�݀��C�ozNF�6�9��A�4�s'b�t�{��7ь
>qob@b#:>�;���9�dՂ���a�+�D�+xX�+���C<I���� %7.q�a�����yf�bM|�GW
_Bcs��S%�];��o3�P�7�x~nG������FN��H��&�c+�/߼��\%�	�zL�N�מ1��W�����I����R'�V AҞs-����H�\^�p�TBG��wx�|Iqp��p)�|{�)�!+XX�|à�Th���*��e�Ә��]�tJ#��I���Ǿ�@3}�j�:�.�O!�d�F ��93�E��6'y�� u�����z;l$�4����?���g� K��hPj'ÅfI�v����9��x���)}�Y���'1iW���.HjFmwƂ�5̣6���Y������t�{�ˀ���;��2�s~�eu�Z�G:S��Z�M�	��ŨD��b75��*�r�%۱�e4� �8"�)v�/���Lk����|���=?���ĉ8�#� ��2C��p$)oY�#�^��{+�k�<mu �кU�浴	d�������6�����
ɑ�`��*�)īӻ���gq .;�竉��4����8[�����Kk���3(��\�gU2ZA�*�]o�n�ʮL �
.�6M�tL�RDn?�6�S"�A��[fȬm2�c1B��s��Um`��d���n��!�D���Z�ʄ�A8s�;��^��Dt�Ks�x�g9�5�Ә'ZU���h�g�l��J�݀���&�UsUS5˳��9 *�U��,E��j툭���
49��!0`�h�*�4����tޭ>�^��ӗ�p�t�� ��o�ƣ����M�]%�T�����<��&�xx��ki�R7`��w#�I��Cso���A`U����h&�P׽�
��F������,/ms����$�@���I�8��>^���AL��/�pp��F9��%��Ane)�9\!'����LSݜ(,��ta��j�,��a��tS7.�weRK�߹TӐGwu2ր�<V�m��wB?���B���3�[���Dw�y�J;�D��p����P�����%�'cF}(y��n+��5̀�r�v!7W^b����'�N	�+��V�����dv��qH�Xbiʖh��o�e�C��:_ ዴn9��L�8-�8ճ�b�e�M?Uy�l`�� �9)C������Zu��k�i9� {�#}e��`���Hu4j��+s��C�D�!���(La�j �X��w<�XlH����O`}u��+���ŒH��ḵ�T� �'���3�/��I/^x��f,4�"E�L[U�>�HG]��#oX��&8���J|�4���^9�j�e�Z���]?����g���#����>��bAH$�JJ��Q��1�qV������[���h�ԫ�<%0���� 3��֎CWp�����ݧ\i��L�zS���q�>&��e��T7�LZ�������Oc�)�з�BQU�kya���,=���\��^�3�z����o��n!���x������O��90P��_�Lڹ`Ȍ0X�V��ȏp>[��c5E&���)+A�/�@U�Ơ|_��]�E��E�v����Ebt����՛��n���P��N	��)���/9Ú۵Y���j����@£���*"�r��Z�J�)�@�O*q�u�1�)u��g�a6W Z��0�/����E��6.L�[�y3O/��FrZ��T;��
6A��ȷl�#t���﫿O��hk��Qf�!i^hO��Nu���W�7O	q_�� �;\�W�6�����>���(n+�M?.5�m��H�
�}mo�u��B�Sj��j�&���E
��,m;����sܹuIb�0wf4��-�bK0��s�'Ӹ��K]e]�?w�N��Pj&�]���¤9_Ԣ�]R8��^�k��{�� _K��(|+#I=�l
,�g
�L/E+^�O�ڏx���6`G�o���Q��(�XЧ�*���fXy�Ͱ��l���0`V�P̰�_������%�u�x�5�G��8(�����Eyto�d#����޺�����1�q�`
�S6/���t���i.D�e�K�q�D����|���<VUɅ�"=P���N���\��	����%g�
խ>G�QO7^���Iу@!��r�C9Ͱ�\|�hOw���:���a���Gv/�3I}��pq��z�d��8T"���Wx�߬�pk5і��q���f��7�f�u�Q
^�����C��F7wz��w.���f����b�3ͬx_~	2�W��ӂ����=fE�Gf�3�r_��!Q�AX>zk0sgm[`!�R�!Uz�XжN\�_{�6k�L������pd0JN�Z�d���\o��SA{j�� �B��7�,f��̪Pǯ��� F�Qm�ӱ>2�;�����=A�dn!Eu 8�U@�-M'�ÿ�'�X�57�(C�=�9�	��rQ�ߤ7s9�.}2\-~�^
8*�k��Z�4��^�%�,$�7][�����Rm��Q�#0&�*D���������^��^�A��ŷ�LJfo��uq�NG~�6_kA�����ޗá��_���ҶgWv��yY����cT)ulΥ���a0'"���IFv=ZdjV�.w�JP�a�׶Aio�})XS�U�M����9U�'�o��<�g�����bo�� �;)����uZ� !��������Y@��3��GF�?R$�:�rΔ�Y��MI�Iw���w��E�S�d�I�GN�J(4(��9�tc���7QΖ�2a�᜞�Y���Y��&�
y����A��l�+Iu�up
�J���k9vH}7��?0����	5�dc�1�T�Kp�i@o��u�ޞ�2��x������#N��,R��y��]֜�6ed�E*|rG`������f #ҽ|��A`Z/��{9e�3�&@̈�  x�T�q��$;1G�R�+0a��H��@��Y�r�w�.QM������e�ʱ��{���������@�dLN�RJjP���}����\�Ff=t�ٙJBQ+����n���'i���uH��"���S�Jψ�d��i�����,O�\�l�S
 Z�h�ˊ����CClǕ�!g+�cs�c7�UpW�Y .�b�?{a z�NA6� >��H�l:�p�?u���w��L���Z��>j�:�=��Y�T��.�\[��I$
��D�w�x��=�pE�ݯ��X�y�=�������\N7U (n��!U� DjSo���XX/���~�K��6�wW5����C�*�_��P�]%V��B�DP(��3\�G���E���_II�N�Om�F��wX�����=j����S���4�����EK=�U��8�N�L��v�$��9H�AX��#Blj�	��ҭ(Ft���~9�񗫆@~TGѪ8��-�Ȕ䑴�zI^a� +T�K�g�e?f�4J)ڱa}�y	�ر�B�֌(Bk�U��'�ix쒙���C�b,4?���Б� }ÿ�i��Q�I2�� m����!}��lM,~�)a���Bż[S���U��fY�rUi=�qEc��*�wU�*�I?(]��*��t5攩�!g����^�c��_���ό��w�\��\4��V�;�Mn�^��>�.���NOh=��o��\�	:��d�pDŊzہA"�H�VT�p�9z�N��7���Z���'�461����nt��6699�S@��_I�]z�a��w��Ƀ�d��y:�t	&J��j�3r'�[~��H��0~XJ��Qy^�O���k��h��i_:r2��3���<9��u�#H���]L�&�����Y�֩�����k����I}$ �	U�6�:ކX�iˊ`�^�2�f��b�X���~��{���v~���z�7$Ů;�=����hM�[�kIk9�O]������/3�����tGU͉�Qi�^,��`�#d6�n `�|��xi&s����B��t�Hڝ
P��8�+s1s|Z,�!�U�v�5$:n�"{e��2�A/�\xm�G�Ѧ��8��X"�7�PZ��ͤWy��d�>�n�,@.Ub�oM���@��j @���Tf7W4<jnW'���~F����}\/�����g :�:3�rA]�%.�z ޔ,�&�%���`���K���\c	�9�T3�v���!5B��'�;��1B�'��'�۾_�G+�7�h��tʶ3\C|p'_��9�:QTUa�Y(N�����]/�?��GNY�� ��!�z �~u���ˆIO��:�8�hm]����tèC�~9��>?�l�y���Je}��8L�jp��Y�絉���n&Ο�]���k9���
e��z�o?n�F��2 ��'��,��>5�!h���M@�(��*h	ő 

�ӗ�F���"�܍qn�ڎ�ҫoOuQo���Hr�k�y<�Φ���~*G��n��I	O�.�����M���h�6
7͂&[^LN���[��C�Ou�?�@;ǖw�~E�:���d�У��1R�`��:n"�p�NL����uN��<'5L�2�Ї�:�����Mɱ�y'o]O5$gV!M{���C�KP�v�ֿ��C
Ҏ������^6�ޒPT��	x�G`�ϩ�
�Q'v-h���d嶁k�F �z�݂�b����5Y�%���,�1m�]�gB�K٧��,�bk؈Cs�jDJ���>�P!��G,I)����z2)�Q��]����_ 2�]ߖ���>��Y��-�{d���Edk���{���Fʔ��U��ˋz�y�`��f������=����`ybY\+~�� {�\��D&��2s��ʀ�@�� 1�*��ݠ�%T�w\����hz�Q���~Ytm�p��D���j��y�2}�tʺ���R��v���ƚ��P�J�Ta��4XP���)Q����@B��+R�F�.F�[�0N�ʈ0�����5�H�M�V<�D�8���MX2�m�1QqL.J����x@�(�-�l5n�����
-��gõOX˺G>����=�$��w�/��w���4����B��(5��q8?d�" Q\X�G�c��^��|p�����uY{EcK��$@�X���>���&��@~tw偙{��B��M�n(���+r7k�ƃ�7����`��xK"�DW����$ns��[�R��HȞ�Z9h��8NZ�E.� x³N����͊�
i.[3�JE_�9���bE���-K��8�~@k�Ŷ�m�SԞ��H��Le��΁����e��h�M�
�m�,�e�*l۱,�Ѽ*�+�����ベP���t��p2i�X��Y�1`}�Y�S �?�%�#�;؎,���sff�1;�u���K$�����Qp�\�����p�Ǌ52'O��<��+�䳒`T����g$/�Z&�W1��䝕��|�D�?�}<�~U �@}���{����y@#���L�)k����*�cI�+�j+�MAm�ܨm���rB�JLȺ-��hT�1��Ⱥ��l�(�#�7/�q�e�8��^�/ڍ"?��[ֆZ5VI��P@^���*�x�Ƿ��=���`�8�٬֧�Nt*�)��%�T�����jmڙZtڍ�,�|��O��rZ�M�1�T�屬i|( +12�-bѕhi����n���nAR?�S�ک�D(�S�T*>B��Q�,O�2��B�:W�9s���A(R�e�}�Wm��_[��ƍ��1q��⻽�0`[�C�%|�_�9��=	�t��^ww������&$�/t���:01TlS���j����,��^�+E\��U6��N��M�=z²,��{ץ�)<|;��KͭZs����	�d�K��5�yĀ��GP@K�p�g껽W�w�@�hsGs�/����	E�K�Z��0�KC�pF!��qӑ�t/OԔ��#Q�3U+)�y��H0 �ztB���*��ˈ?Ʋ�k�n=�)�����ʓO2F��F����-66@��J���/�����D����0�-y�O�������X��@�]���n>�L�"hڸ(����:f������3D�h�ϐL�G�ވ��@�{y�!DJ�q'�F}�b��4
~[N��i����M;- =<���]���o�ӣ^*a����U�����vЀx�����+6���n����X��gCiq1��C&�4���M��jԁ��;�_ow�G�z�]:I#i�I���hD	Ë�������<V��	�Zg���u�Y�MV�Z��	1��e�7/��{�G%0����8G����xJ'�*Bo���x�W�9�`�%����䏁��v�Me���`D�,��o�k&���"��z9�L�����&��#�Y󣽺��	���0��ډ�����L���ϣ���$�0���(γQ38<2���Sk�N/�h�cVeZ���:֧1T���'�fm#��<�͡y8Ph~JWL����̶��c2�^?�t����i���>橆�+���?����׬5���kl��pr�o�t�������0+���ܵ���K����N!}%1��9M��zO6q��/�N��;�iѹ�	�Ó�",��˄#����S���K��g5��a�[��HÃ�#ٞu����n�\���٬�AZ0��*�� �@��e��+��y�zL{! vލ�7̖c� D��-�譽�t���$gUh�@ܨ���	�r= S�ζ8I�9��TITTe�M����Q����Q��렅�RN��趛��ҷ�:m��C^0����ID��2���{cEP�_4Eϼ��"�&�ِ�e�Yh�<B�7Ԑ_�V�I+���5�_�B�n���:��9��N7n(e䕟�H6�?u���h%����m�:�RP��H�t�Q�ş�<����%q��d��W����Rx.��u�c4�@��9C��{�7ԁ/<�54�lC��/P�|4��	�0(�SS����и^��N�v9o-�L���7��6kG��M����%�|�y:� ,3V�6�@r�ſy�B֏�E�Y�t��o*Uo�j˛�so�	]9n�
�aj��P�k��K������I��ke�cE�e��#�7�~�f��T.���T�뚼͹�r`y:Jަ��/�&���ڝլ�8���1u0�o��� J�%�%^�e�+dF��U���g�æ��Uéİ�ęW��qM�@��|��ކ�1�P�d��w/�� քc�Z@��������7A��r�%~N٠!���QuΣ{}���apn�y�����bdp�u�:��}��u`��T'1������A�Efw��� ��=��3S;��aV��H*_�Ώ���ui]d�g�`��"G���RI��2+��/ؽՈ~��E��a��/�i{�����G&@D�*ӣ�!{M_����	����d@�������>|���3�M�p�c_6D�p���<���5�Z+}L�Hҽ��p�Ǣ#d�%f���I^�p��ە(nL��sW�Vf~���������l~�9�6��;��qQYMmY���6�̼F$�6�q��������������ƛ����zh&T:�X��*��A�9(ؒ�����'vP����WhNtB��I2D�W�;��+X�'܍��K�UF��#�H��F�
�s��w�X05 ��Ji��l���ݾ�%dS0�.`|8d��1���u/�Ը�Ӳ���n�q��SẈ眩��X|%G��\.!�w�$���XF��3����%y�£���3�t^�Ie�<��'���0������0�ń�BEDvw��]����q���c��:�:G��AP6�fS�
[�S���E�R��1���5#�� v�K���+�S蔖�y;v�XI�1\K�7u' �=�(,�;�-���
�X���=�9ۚh֘����,����E��	K��A���p%����;R����L�>1i̉}��0�x�h@Q���iE眕��*@a��q���!U�3�gf�'4s�Vr;���wZ��TzB]�s�P�6��|( ��	 ���G9� Q镵;-��oQC�$�\�msFMh�} m�ɹ�G򣆁U�VW��	)�b�awT������';]�ʗ�C &S4C�:E���^tI�קZD�S�����䬰%$����ű�I��������	�v��ٻU����Hlk�����V1�^��e!��/��ԏ��S�>M>j��f#\��K�d��˫1�ɂT���( �=��9��s��uH��'t:by�]�o�i\N�sk�v�"=��ǏiP�݆M���;�[��Ò����#����g9�KO7����lo��4k+�l�)����UE������-����%�ztlN�s�־"��Fv�6�ڍ�TW�ˮH�?P����l{x{�v5ܵ*(�;wy�^��|qu�U6��*br�H$�RY�JC���%���v�NY�d���:�b9@�#gH�Zj�V�4� M���xv��f���z�A�"YMD�#p���5�VT[}[���$-p��L%q!�$���y��4T?qݽ�d��~�R��Őf�_UӚ�m�)9Sc�%��"�q����M[XwޢE:,�Nb���`��CP�X�.-�e��nѩՒ��\s�;��6�g_�	���Y�j�L�&�d@7�R�@U�sl|8��b����Y5���<)��c~�fh�
JC��*vç!�Q�gk�n5D�7�D�$�/0㊋�)�]�OA9A��3���?������o�Sn�%��P�RoL]JVX��,�ZQ�#�X��{��ߘ�T����-.�cz��6�8�-�K6���Y0��i�,Ϲ��7G� ��?u���)��nw�7��ͫM��#�h4o��_� �q~�Ƿ����a9m4��(AM��j�c��
hӪ�dH�IZm;��Fz��lh�g�H��Ѡ�Hq��hc4Y�6*X�o"��J�%0tW�.�0�-_�qg�����vA#�y��崜�7�b�Џ�	T��^X\+T���c8��>�������	�pAS/Jz)~W`�[E����*���w�xv����EB�}�Ǉ^�i��v� ���\ �w��� cR�ږ���F��
<h���}g�[���4Q��G���;���J��*'�X#s�3<�7�Y����I��rv`I�˲���z�`ti�
�=����
��T�2����[���h��T�T��}��I��y熪�Q����~F`�~ODlB�s`=���[orr��c	X����Q�7�(��ɡ:|I9j@�y;|Ë�7���9�o�KY!:jKe
�5�r���U��ҋ��dk7�F':+!D�Q|3ԁ���!�H?[o����M���6p�5�����"U��۸21iS6��W�����|�p-0t�o�tPyx�:�{�2���&J��X��2���wf��)FV�Z4��F%]��RBZ�ֲ�u���B��6�7ן�萓�am�D.��*}�����Q��{���F`"��t�肓��`�3ǹZ�m�?�M���Z�pi��-�mb�dr
#dKX�-$F�¤��e�/��	��o�/�:i(����:�4�JÜk�@�5��H�e+�ptc�Ϥ]j{�Z������D�X�m��=�p��rL��cx�{�띪*	D����[��S �7K�^0��P�o��HNc{7��0p���] Y��v��Ī�m�!lxOTI(J�p��S?`�FV�9I��]�Dt�K[��Зq'��c�p��� �f��!>y��f4~n_�6�Y�8�\�W�,��HO�A���U.��6��nErav��M�jh?��G�y+��(;�4��&�\:��`f�i"J�>��˭��y��s�eo���u�����([��ǰ�U�6�E��&Kʟ�:%5Yz��a���bkiNᯘj�j�J�3��P�K�9�9�bPvi�z�����T�R\W��)��:<���I3���dZ�Ny�7���l��瓰ޕ#��m��^��>>���p���M|����z�o��	����������:��b��H6�Wo_�"��k�vy���4�=�����?u��	���aO���)xx4(���U�9)���l2�$�D�eo\�;���h�|v��_ɴ_4����>��q(�J���A�_i�����x�J�}uy�ś��՘����,r'�.�塒J��8<}��oQѽ�����j�+.��l����:�u?�uX�}-����U�Z���8��r�V�j�ω��O��1��N����G�AU��A�z
�G����ue'��_�0���ء!�`����x�����Y_�\�x���93��$0��! �����wMW1[����x�IDPlI T������蔉�Ѝ;W�Xg������>�Շ�6K}lߥW뉟���z[b�������Q^�9}52�����k&�w���橍��m�u��*�!�HiyC��M�p�M{=��Dj�⩵��u�&�X���]���rn���2�* NDk��Yr�YҥD���1T!�/�v`����Jwyß�����\�y@,aUt���f4\jL~��!�8���.\��ҹ�ֽ[`���s�d�Aa�l�|��Cp[Ⱦ�q��^2��^�8��,"�u��LV��/e׷W�`��Y(a�q���.��uú_F�U�˝�X7��Rۓ:!b(��HA62P��tFطIm4��L�F�)�:�3ڛS#� R�[q�������I|��mY�G�%W�pG���A��6��!R��g�s���R�V�g���|-����������'Wfj8�~��:���f�
�ԣ����*���9���tHH��	Ŋ�!��92ڹ��!�q-���;�>\L讘B�/n���-"Z�nj����w������X�&r���`n�PLُ��w!�=:`*	M���I��|��n�Nha�S�~���*=�T���Vudk��N��� ���{f��w�)�g���/K�/}*�q�U����ѷ��!i\��$���0�uɀ0rn��`��<m�#�	k�1�D���r�>��㸷��p�y
~hs/�w{�M�-��BFQ̿�S+@[Bcx��T�g؄+�ѐ�����k�ȝj4۲}�f|l������<q�+6S����\��#��D�E�A���u^{����I���4Ld�v4G%+�O���a�%��i$��pI������1�y��# � ���h?"�ZO<���g����\.@��b��Rku�bR��~.J[�#�>�<��A����s8I,�&|���(�}{��RR!G%�_�y��i�.�,��t��{�5����E���m���-+�`]"Q��!B�ε�L{dd��yP_�/#��t�J��5
�g����,�8��?\ކ^*7����ۣ֑"�#:��Za�{�H�+�2Q'��8&�\ƞͻ��8cp�qp�'�L��@п�K��5f��u�O0�&jwS�Ͱ�d
w9�T��dY,���ֹm��R�O��z�!��RP�/�N��*^۽�N������k�E����Y2���e��].�
�W
��I��j�7`i�F��hG��d��'���]x�!n$[�~�2s��]�M�w ���Q��״Q~n�T���V���e�㲷���1��*�5�3M��VPgM )�!��K�,}_��]�s&/����ȇ}�S���.;ᓎn���K��E;k4&-<'���J�k,D����baT_�Q9��7��Y(H�ĕ(kw���˖h
sIom��a��oz������pHÇ�mɯ�����`�&P/iߢ��w���'�2���L�?�HXsր,��U�	=��3�S�x�0��.�?ג��J0%��-�������{an4~�K)1��3�/��TP�\n+�
Y��5���_�������z+y��� ����ukǙV���`�̨S'���Xx�B����wދ�v߄��wr%v�����i#��*<篑֣}/Ğĳƺ�Lt�d�9��7�\��2S;��)t�IųuC��g��F��<�&w�w��f��E��P�z 3\��¦�P��P��3列{�S�:�nn�O�ݐ�\� �ԇ������o�S��B4 ���Gf�<DMex���UV� ����>6�K�~�A0 �<�^�/��_M��v/�������>�����6{跰�j�?U�ȏa6zy'Q@0_&�C�C��%��X��3�����/�uA�A]�对�`h�ȡ�>�`p.�π�XK�@N��^*�?�	�^-�
�l1.���>�yK����x^�^z��^&��+$߶�a*p�87���J�T�<�]����\�v$g�-(Jt�i��巘υ����l���H�����	N�w�A���UЂ�8{	CVs�=C�����l?��!�7]���Ĥ�C���)��K��~"g'�B(~n樂\';�S�"R���њgTDc�r��u��8����!et�趹k���C&E��@��f�$h��r�Ɯ/>/U�u����G��)i�N���!�����{��v�A����-�VR�SQ��"�}�?��S㰞����m��4�����~�V��3@R#�1%@��L�b���e�������I.��i;l-=�XR,�}���0�{��8��`���NՒ`](�v%�!����5y�&��/>JC��y��.A;�N�/�'G�&:��r�&Ko(�rjS�hA�j�[`�Z��O
�B{�QЖ]� [�?&+˸�p�-v���g2���4��:A��.�A�#O����+�$�X^�g��� ��4�� �5+�%d샰��HH�Vz�8+=�>�%d;s���Y�S'���f5إ�-M���ׄ�yA�~t�	�)
���a3}�T�����i1�d��\??�����s�Ζ}Bp��E��\��W���Jf0�$���[�a�ϠTuO2�[�A�eù�=%�Lix�<�@$Z�μ�a�����E����d�������Ψ�5E�j~
�<���s�F�S^�ݓF �+����4�7ѯ�\���R�����C���,�e����d��CbA��67?�꒩��f��Sۉ^q�B4�ʗPcج�J�-��,��!/��d�^�9�e�g�!JOb���RQ6> �sacU�!��W�hʡf"�Q���LQ�4(�F*L�e�'�Pܒ����Z��[��eE��?�"�<F����f˨&�Ϗ��G���������񅪯=��<���\v��I�]��gW��;�&����&骟����R)�����Qw`se����R�N�H3-&~m)G�����Su�Sǁ �m�MG���S$�<���	�����<��9a���a�n + �rxB�7��,`)Td�>7���N����B������:7����'���_ޖ"�y�|��z�8ߋs���k^�N_��7����łb�.�v�$�"�6�-�y,�E̿H��Y�@�7Y���O��d���#�!��)��.U�O���R@�gE8f��@l�-b�2�=�G7�xq�k��zY`DǾj��̽��'t�nSD�$�3T�W
�$6�C�K�-i���a�]Wb����n����g@7)R�A*ME��;����F��U~�������IHS�iLT���h��ի��D" �s��r��2<!p�(���O� q��2�g�ބ��ѡ�kh����}Vg��M�F�L����B��Uj��_�%��Ӈq�=��F����8���-�V�Թ6@�D�F�&W�څ8�r�@�5"!�<
��k_�����/'�<(��a�:l.�iӄa+�lzi_.@J7�_��Ɉ�~�$�׉����QJۗ�ؐ�G�b�=-{�ڀ0���H-I�7��D�ޤ�E�^9*�#���( v=��M���V�"|:._�N�6���?#�!s'�b�:3�H�xe>'k�[$���&�����1Rc��j�wS<��JQu�w����EZ�m�Z��R�D��f���b؂��t��F�5	���Qb�,����i���}Y"p��7@fV�W��Qq�����yfJ.�"_f8NrNRM9}����鋠�Vqh��]�ܔl+�7M�ZM!�Kv���l��;fyL^L<0L�6�P�+�b+��x�Cࠗ�DOSf�Vx�k!�>;V��V�2q]�sr%XZ[e�E�:u�6���|��#��b�p9!�(U�F�c�n]�@|j��ǎL��ӄt }�(�$��	B��6WT��wY��^�}���\�ԫ�[���%��̚4�"�m�Q6B��Tfn��,�je�nG�*̗�*(���iȕ�*�80�+�Y� �=O(��n�_�@1Τ�q�t�h��A|��f��:�+�mt�2��ƇM�������b}�,��ٍ����/��s��*|�n���w��OIY���d^�����4��Ũ	��q�V����.�-��$�\����_�oBC���y��&xT� �G~�⮥bn�T�̛$�����Z�]ᠰ����)�c���g����⍱r�b�k���uZ�����*!أ�����wx��nnP�c���G�?��w��?&��y�:�Hh�C+� [�����Ę$ɵ�B�-�-B/_����Og�Ш������[�.ex!����1�>��eD�;��K���jF�@%OC�S4`V�����]ad~�bU:+y����)f}�DU���s���	���� ��J>�e	X��G'�8|`�����7�.4ܪu���=Q�"�c�%����f�����&	��:x��{2��ň9�lJg�m\�od(��lBij�m�ڥ��}������`�/4aܢ���=Q�W@�J*�ʢ�D���E2��o�D�4���?�J3�6>�	�wNZ�FVAˏ�~-H"���"I̨˫�k[F:u�KaJ0�5���J�Jh�����}h�Ew�h�%S��FS�K$@r�%�m������tkN&��r��:�6�eszU�%J�ՆP�xl�ٹh$=��L��S��P�P��^�z��~U�tɐS67xE��73��p9Ȋ�Eg�L˕�8���˲�pL!�n+�5�(c�焠�G*%O�=
��j���I4�����<�y���Q�M���߰D?�ε����Z�pl2������� q�~����U�ۧMK�Jb����x6�!(�� 8E(I�#���2��^�j+e�7�<"V��Y��T��(IQ���a����$�*���e�kK����[���:9�y��a�Om%�DP��؂uhjv�-rte�lIn�+{0`�^�-���<�q�~�ߘ<1�Зo�jY5�sD��-hوy�Z���Nc������Ƹ����-�m�
�pS��\��8Ѕ��t�N/8e�س&ۦ�ʽ�Ҵ_Gp���x�"'�/����-2!0TB�]�:�v�.�4�<�!륖Em����x:4̱7)d`��y����E��<���xd�Va/��E`���}��n��x�� �
�n��o��l�FϰI���@S2�zE����1!7�j	9c^�'�_��3#����7����&�rV�׭�s?B���s�+׎�	�ڄ�a�CE-V��W#��<qB��.#@X�F���]�g8w�V!��D�~yz�S��V̴LN0����j'��3�4n@Nl�.�n��9����4xr�$����[m�x��k�ש��x�V��°'6�GV:2���bb��QHC���h
xS�!6T����k�&_/�K������v�dUȗA]�/Qv��`,Ĭz}�`���G�жB��)�"�f�$�����*RXM���:�SI�;su��KQZs��>�K��[>���a�٦�O^Qos��
ei} �j(��.v�4���61��B�$��Sg�����MȤy� �i�8ܣ�1��p����n���S�P�T$M���rվ����2.S,�ssT}�)���F�zad�������?R���2�)r�K�F&�g�޵5��f^�?7��Y�;���'�J�w�u��h�V�3[���7۸`x�����1�����u՝��@� !���	"0DMݹ��ff��^��D�a;�i��(M���c߃S��7�M��π%��Y�����L�C1�G�/=��n�>�"����e�������o�eR�j8s݌�21 8��q;)�2o�5=[��v"�%�+�3�K��_��el��O���<�Ĺ���
�Ĺ
��##���~�U��E\f�n�]_j�$�u�݄�v,���K�N�ZbG�0��t�&��i�z,;�)طS���^��~���Nl��L���[����I����붽�.K8�Τ�k��,�h AO�QxBa���9a�,�%?�P���mֶ��]O���qZa�/Lv��\����=RG��>Z 4u�$4.��{(�Pl�`�Y�W�5��r!l&�(����ھm�5��d��s�Sosc	�s������{8�!����C,�>����x�QJY��j�J2�ab蘝N��2�y�6���q���,~O�xO��7�7���c~3�c��g��e�*�>lS�����;10�YK�����\�ל8�R�bvD��ٸC=:���?̜���$�!��1	��ӌ?���$��z����� Wl�e��,X�7=ϓ#/ǃ�����|�&<�*���+\�5F%�L�f�m�p�����4�3X��9FPJ�d��Ȁ?��P���1�� K��9e�σ�lڹ�x� T�Ή�����/p_ou��r���V`(�Ɋf�x�1��r��0�N�JB��'v���ʒ��Q?>���y�M�غ�A����ܱ�v_Y��
E4���WxԱ�ku�b����)�d��,9|i���7�<���+��޵+���x� 2���%;�Rc�%��z�K�����4CF��E�����V릞{MJ8L�f5`z��4���C�S
P��0.߲�R<���� z9��2xxz;��+�%�����as�ƍ͟Ϫ�n'�����%6�{�eZ�=����v�#�}�GX|��{���[7Lz�ł�䧬�3��4߳
d���1p�8����@�lS]�w�,u�o����gQuqo��������A����>��G�k�)"z}�Qh��$r> Hɕ�?^�-5gO����0�l�7�ڣכJvDv[N��K���4543��c���[�p�-�ou�������TLb��;B��΍MA�e�Y��ǌ�<���& I$ʯ����K�[���(C�?�l�d؆�tA}���طgr�K ���h���>�Wҍ>k�4Y����m�����E�6�F?���Z���������Vm�xt��p�p��8�p�m��3�ސc\��T��G,R��#��!��c��4��fY�ӬZ�zDJ�.5;׍4#~���Ԭ&��J	R��NM����/F���(>H���@JZ7�0�&_4�71�֎���-)��{%?���ߥ��q�^=�Щ�T*��������%��'�
_�~�������%Ip�|��j?!�7���|L5_{~ǂG*�HG�ˈ���>Tj���O־��S�笒����
�@�(��ާl�&�3u
Q ט��i:q��9oٹ��)��Kw�}����<hD���>�$i
�x�L�����L��Hgz^�z׮��{����ie��
j�^�hfqO���m1շ&�@
{��vA����[��H� �s���z,԰����D'���Ad��d�x�gr�A�����ťL�s\b����l����O�oϤ������k�;�0\[�+�k�H0��k9n�מ�CQ=�5��v^������&�E�AOf�Gd��P���?��Ԅ����ϭ���ȝ��a����k'd�W�3�#�*�G�4�.�� �kX�2YEW�I�➳�-�U�\�����&&|�ي�� ȁ`�����v)%���Z���*���^�7�yã����NkKY��
�}��w����ZX$:��9��a>�M;_�ޤ�����p
^��]ʙU�堈i�pdwz4"��I��p�%3am����,&u.Zp����L� t��t��N����\�e�S`��?�RD$���֥�ַ*M��_�:��S��p����Ŏ�'��-�h۸*Ȕ�Z�ȋ*��p�k���j���pN^�$�X��B��b��Ob�]���S{�z�!P�YPmH	�:�%�z)�ɕ,�Q㜌��Q�X4
\-����B�R�ļ7�3ace�&Z�h�@Q���?�G��I�"Z\g(8�K���P�Y}:����|��/���N�ލ�_�{Ɣ���ͫm���U5�
p���;����_'�����,�95�Y˱n@��!��76�~��=���#@W!��`��B�\9���>{�e��mA�����*7�BŇրh5��C�������f��O����u�u?��9Î��{{������d�yZi��U�Hj�dDK�<���oZ�ߧ���C�=���Y[(�~��:�?� =�-M��?�P'�n���5�I,My�����2�d�;��#1��{;��06�] �%�� փBt����~����[r�	�F�!����6�[N��	��)M��nW0o�r|�N�z7,��&���ʽG�PiY��wd��&.�[t뛊/^�	��-�0��n��v|�9�c�)mǖ�tG�jv�+��\�2�Ĭ��zB\3۵_R��)nn'g:t<�u1+���҇�k6"-Uf��N�ri1oG:3����n`�&�j�	`h��cN�^�0\�m�	��s.� 4tP08>��(�.N�o�WZEX:���D�L�ʂ�¬n�x�(����2{fC_[#?�Fn�,W;�l�/������\�I��~&Yh���_G���{��!����Ex�qގ)��D�?�Y��w�p��*�x�k1�i$�i��``�̩����Y�ьn���[�X���eŋ��hu�3�&�uv7������P߀Xӝ��b�p�����4a�I�0�t���s}W�3�WgM��V�X&!��1�.p;sw=�;�0�i%�)Q)#��}v��y��G$�Js��"w����}�h�$��V�.0�ǹ�0�;�R ��8�b���$՘]]l���3m�Y��A����AD ��z�ُ:�$�lj��,'?�F�!����m��͌~Q��r���rV��r�F��T@��F�����G��>yk�y�LA��
k)�b3~�"��2w��ʀ��]�Lly)����Q5���ĩ΀�Lh�˟-��檂
Duږd���$6�� E��/�)���(-��D4��E%[s��[M�"�J�y�0�~!�������ܡW?��͆���$!�6�������d�ϕD)�t�I����w㞮9�j�ߍR뮋����4�è����vc�D����~�hu��A���w"�^�lo��L~_r6|0�i7��H��D�t�\�A)S`��ځ����Xj�im����݈�3��t<�j�5�4 �h	[�c<�%f1Wބ���ȏ��(�=�A��_ 
�7.]ZM&�cl���X�neٛ@'(l$�+�i����WN�y�MP�G��Yߏb|H�+���n�����qɳD�����t�X�m�B�d�\H�c�� ���~<����m�C���G{D{B�Z�,];�iNgL���M�|_�d�HZѨ87k���ə$J�{zטo�}���Wԣ�yL�lDa���b鈎�=�jIZa �D F���StG��Dz��55�iz�F�dWq�(�,�Ek�@-_�)�^A�*@� O���Sxt;kd �]�wN�$l�~�!��e>-}�@5���ꦬ�A~����H
��Ӫ[T����������x9�	9Ⱥ�c�3�]�R���D�%�����L�3]�O����G��O����<�s�֣��ք����c�K~�X[�v�@놁���Ѷ����4�:b-�|"�x�z�d�n.oy�����̺�9����b���D�5�Q�{�YѤPކ�,ƟDGk�+�%'sc���A5&�E��n{ �P�߫��ӕ��Pq��-y�	:���)�?N��)��W�~�7p-Uk����lx�'�/H�0?(��k���j��!�IM�I��r�IΐZ^�`/+*h֩_|������$���(��`� 3���Y�XD��U�����x�0Y���h*��u�D��bIb	�&�]�m,@��r�#����a J�x�|GӣH�+�s�MQq_��B�����;±}��(��sW���g������l�ZO�('��Q�������{�U$�T��o�_�<zg/��klfdo �������P6#K���:{MU�/ ��s,-�#��[�0�ˏM����@�`��K��Ḡ�'uS�Dc�S�g���iޠ��_賭��)����� 8ݺfl����|rbQ���D��řƬ���Ed�Jӿ�8xa$-fK�[G���w�� �;�@�^)�~D�,7ڧf޲�iG�[�a"��]�mtYSK�o��=qǫ�0#dg����L����c�^�\�'�|�F#�ѻ&�B<���I���ؗ����+�5�Q�8`$R�+hGT�-�B�&���3(�{*�Jna��Z�@Kg�a?f���q\b�uqIܗ1,�G�K����g�-�i	tQZf=V��ָ�Sn�!e�e�3��ӎA���;���2` Mα ��f�C���,�Y�VA���!���%����W#:�Z1˴�a���k���7��Q�&��LȦ��`݌��i=�,bS�f5�٘ئ�ע�։��ʀG�R#��wT{alƙ��,��Z�y�JΚᄣ����9M�2��a5������'��LP��S��k�}�_x,��)�D���|8�����%"w��\�}m����1�S�2($��C	p�b����o2���:.$�tm7�O��u��&�$J��E�b�.�P�MN���F�fM
��g��Q�s�7���	�aO�7��"k_�=�H黼F�$�W����������H��)R+�X�?��N8f�Vԯ�H@˯>��������%��%0>3Ϡ%(�<V7^L�Z�馉�^���}���\&֞\%�#��D�+D�K�WC�lQ��I�G�� ��?��1 �c�ҙcԦ��;�u����Mj��i��0��(���	b] ��#�I��Kɂk筩�)�����"a�֖&���7�g��@o�	ܳ�j[��"޼��,+u�r�CG�D%KWZ�8Q����DӮy�n6S���YE���eQ�"϶�m�E�bFHG$t[�}ҕ� cґ�H9���G�ϳɻ>~�O"��(W�#?����P���1�t��An�'  ���P�̋nX8�<���+H�����L?�?�⁺�v��h���ʹ�o��� ��R��f:�˧�cF�r����qW��� ��j�@Bm{'��v�x�Pҋ!��%9����=�Qv��{թ/�UXd'd~��r�׎f���*��D�1R��}b �-퐸XV��D��Sh=TV�TkDel��Q�wiU��!/�˴��g@z���y1�����z���c+V��ho�C�2�+U!?*o��b���S��d_�ѥ>k�$&���Ǭ��I����D@����)	�����q�A���{����r���I���lѐ��-R��q���׺_��K ֊J�}�"h�.J�d*\+�=?
�^����9o�F�t�cW�b	lF�9�=��r0ZؓX�J�i��H�B��P#Ye�U��M��˭ˋT91�LB�Hv�m*������`ôЉ�Zt��i�R�l�o�"2��0�U��s���0���L�c~x�(KN³�` M�+�t`��#@�E�1 !s�i�c���)�?�W�R���� �Zλ|+`�f¾Lm5>���n �-��c�n�'5��V_���5���#�7Z�en��$�6���.М|��͝ ��ɴ&-�mR��5|>�bL&^X�Z�����籝�HF�(��\�L�H�?��E���2p��]N)ԁ�
�M��(�m�YT��X�&X����JO	�W/[���i��[����:|l�P.��R"���˯`m�k��xhc���ť�>L��)�������}�V��{.#�	��3�9/�(:�[d�N��.�x��cZ��l)i���=Jw��K.V*C�w�>e��Rgk�%�e\Y���נؠ��Kܢ0�P�}����{�jy������" �]}z��?E��N:�W��<�Fڞ�?��5�{����/7*	9Ք��/�z�w��C�w�e3�S���ٗ�J��k� �[��� ]`/�o�4M�H�]͎{]�;k��s-�����p� jT�U���-���U�����ԢC5�+�zqS�>H��`M�[6�3�w3Q���5<`�����BBWg�6�$�%�aC9��7z+�{��	����0��@����jh{��[M��&������VuS~�[�L��3]R��P|�Y�Q�w��H�cV?�Q�����.ng;�E��ύ@l j�E���F4/�*�
��N�k3K~N�R�55
=�	�yz���s�g� ��n	��N]���859ǖy��7��8Q�`���,�@�>*]�����%���J�40�+Z�PU���]�<���H٣Ⱥ�3Ay]�}���>��\/�Z����rzU$����.�T\� �euǩ�8G���8cj��0��xL�bӬ�m��j� w�j�;"��j6
QZqBGuJ���Yyn����,���������{k�C}��d9pї�U�<~e�x_������!��dQQ�qVu^3*� {��*�F(�My��g\��� �3$��g��!�,��g�}�"&���9�#��Z
�����P��
,׃�*0I��)�3w6�H|.�U�C�,���`�Ŋ8^y����lKT]�Ժ���3$��X�1�ys�ԗ�ˇ�Y>Eӥ3~��{?X�X��Y_�)˝ oK�ꚏV� �Tf�eg�=Q�J+�'ꌣJ4��g@p�;����6�\~
�UĠБ$ ͧm�)�gc��T2���#˾*f3�`vL�Ub�}�V7���?P���E-�u�p&̆Iqc��>C*|�2x� �mt(��/Q[~2�Q��_	.�^V�]�K������y�ly��	�J6��XW��	�~n�8��L����(z_���@Z���䅏���嗰W8�/�|�̕����[F��)�+�
u �]YՠO'�>[���[�T?3&۫{���q>�G0~�ǰ��Z3��B��ZݣL��� C>�Y�f�Q�]�:� ��eQ-S�t3�^I]0�JU��Ι���T
|Jp]z�<�n̢z�3E�P݃������1��ӧ�"�Hs�g��^�d���KN*��/�i��'h��Ȏ��Q�Y��[�'g,����\���Ŭt�
�u��#0
�m
�@���� T����o���|�J�!<�4�8Od��L�w�E�1��ߏ[Vv6�U���շ���>�B׶�jۥ������S=ЇDoO]�C�"���������"?j�O�7|��8U�:���t3�%|F��w�q|V鎝�B�����I�@n7;�Ժ���l��@�����`\*	�&_�41R\]@��s�{�Z��~�%X�;�,x���4.ƚ(�a���
����P%�A�	*0�o�q�����@x}J�^8S� X�����^�QS�)�������%؄�K7)o�uFRn)b,~ec����DK0�O�`�h=��nj�>�0�ꎭ4V��;2fG�F�'��N���:	�����@�:Lm}�ۮ7�pc/OE���'2y�	��6v>�RW|V���Щ�(��y'rn�g���2;�!��2�O;��Yq�ӑ��G�c6�\����N��A����������Jo�Ko����W�:��͡2�}����%n��c�A�a��~p.��)�Y*��zІ=`}�"�`�+�9���X �^��=b�W�)NX��܃���I��w�eM�c�����eJWDqvkY:ܪX�N�v�2�D���{�H~�JFL5+V�(�e+J8�^ّW��Z�c �#�0*���0��aTKը�q����,���iF͑��G�GUW�L��-0O[��������@�
�K�{���S^j�'x���v) ��XE��S9ϓ����u��й��n�Z�Ԇ��׭���&m?j���j	uͨ����D��ݍ�㿩���@~�y��e��}�`O#'�;�G�Q}�@X�:��,~HZ���m��\yO��Ϻ#��NLaD����*�Z$/���W���b��q�塕���� ;T�g�pǊ7����W�R�d�P"�I���5 �]�4�mzIj����:W��p~@��,��>�N��oC���T�p3��/U=O@�ѽم�-�X&�fT�{��G)���`�.��L��ˆn�ɖ�!;"E��X�Ջ�G%��Ӗm/��8H�,��6_� / +����S	��%�;\s�I�ǒ�)6��,�� ;$^;�_�oE㱀D�\�l&��6lm�sy�
�k-��x¿
F{����$��2�����<��ӆ>��H�M�^!9���(�����?��8�I�L$X�1�Q8�4Bm���J���;��U���/�<�@�>��a���Sְ�隸��*�8�"�8�6�b���������!Z�
��!R^�"�Gfb|���20B�����n螌�XGqk��O��B�'XQo�TA�Rdq؆�%\t&PL׾������o��|�3Ex��_a��_��3�	�	,\��:���bD�F�-.�:8�	~f�cZx�N��\(�" �z����<J�[N�{�sZ^����/�QRCBHU�s�D\�h���Q7ʐ?�s&Ewll�����x��ݹJT���gۂ!���ҷ4�!<�"FY����X2v�q��f�~ރN�{Ϗ3ج��^�`Җ�]�l�L7;�9�^֝��|���D��$�]��⹢�`z�OH�S�B�};G��isd׆����G[HN[g�c���UAʹTw}�Tm&��py��bO}�rH�dx+�5��M,����E��l.�w�;�����\w��D����D���';W{���QнW���*T"@�s�M�S�t4�ŶS��&�D47��2��t�P��M�U�;h[�E��2=H|���.Q&=�<��S�Q��ӝX���ߋ3���:9`� 7"h�㹦��6 �~_0+���r��^�o"��U��8�dݚζ�>�Č����8v*�Ÿn�{�w�����ҁ�{fd*�@W 8E�����gJt	���r��`N�O �3�<(���4t�|���`������囔�`P.����s)����c���j��{_3��"@J���j�A�,4v}fZ1�S���*ئ�ǿ�0W���]����38��#,��e��դ�U$� ���Vgd�0e)����-�u���#�w�;ll��)~���L���ؤ�@ ����P�����C��Q����N[8�oU0�B�
��uX�� J�4�������9����ٔ���1�H�Ę2!d��½)�w�ͻ�҂�W�ݐ� ���~F��o5��$�Vg����>S8kכp�9=��{���^QM��$� ��R�N���m(n�.ǚ�����n:^�)|s�O�.�-��Ơʹ���X���/R]��b�Fh�p^fa�.�~d��I�7�s]Vt��\�i�s���5d�&�RCS�)��JFi�ŏ���LM���L,��VpTm����.�Dy��t({�r�n6c�6�*>�`�b��I+�L6,Y�x�E��!�8���zlI��lG��&���a�#�`SUI�k�Y���2	%����J������vD�ָ��B���O�8Dqngg�-O3�:�4�=·�Xw�Sq�%�e�֏�x@Y�]Q����k�'7���`A;eܙU0b\ş&E���Y��)%7��a'!aF����st��P��5�BT��I��?`���Lr}ny��ߞ��@�a�J!��D�V��-���Sk��{Z������*�ˠ����nt�����\�=�'�@�`�-c�2U��xB��34��C����Q sB�%T�x��yᏚF9s��g�>�v��	>&'#iGN#t�
	���DJtԊH��.��_��4�h�}������=��F,�YD	T���K���8[���ut��qj�f{�Sg�%.A2=9��M'���|���6��SZFDY�<��PW�#�҆7���he7%�y��8�xe�_\ �ٻR�5��IUah+&����<�@y?��C�]���׷�B>���������f�̧�?,(�+t~!k8<�%ZwO�Q��o�����'t�f-3R.�[^�U@>�Rap�_b��H@F:���5�~<m𬦘ώz�u�?nEe�7���)�#����>��U���|�ߪs^)���X#M� v<Kt������)��Y&/0ޱ�^�]�a�_��/���_�!e�$é�>�W������ew����5=j���V&X�c�D�.�����Hر�_DH	8�9�|<s�~#Ue�V��j��x���y�CB��V��jV��xL[�.v&���/�5AN�D�~�h��dJ ��;=��Q�� `�
�o�.�w@�@�y�A[�)�mAb����)y?)5����qsc�	��;�[�ؐ�=�Qɍ����'Y��H�4�P�ꢖ��p�%���.�ۍ��/��/�:��G$�j�F^:�5��b
}��u�BF��.���Fu*���|���Hj�J����<�Ż謠��5 ^c�L�=�v.4�S���ZSz�B��dt��[��c^�˙�����n��ѭ��ʊ� ���w��!�5Vx��|��!��� ���Go�~��}�A�b��ZOX���ή���B��1��ȔSfL�!��A��3�EŰ�t�zX5|�c��R�����<�!XB�8���3�F�>��؊�$x���_׿j�P
�Yŉ��Czݏ~Q�T�po#1�%����N��~;I��̕.HcE��NE��S�W١86��A���yZ�ׅ�Y,y&��4u�N��Y����I�p��>�jJllT��ڰd�z��qid%Է-.����<����.N��|T�僈"aX���"���T�o���{����c����j��������N��f1�@9ZEm��ɞ��=����i��VL
�1���UPL��J�d��}�g�b�����=�Y����4!��_[�N0v{s��:=v��)�"���X���;�y������nW�.|���2����*��)ݿ%������5�_�JS��4#�8��lmL�Z�k*F}�*o���2糿�ҳC�1�ڄ'�̦b�-.u٢MA7��r8�
r��x�s���dK~R�i`>��6��K�2l��WG9�{�^��`S��C��U�}~t<��Q��!7��s���Ky0S�0��G2$�hg��D�M~�d�\�ޭ��PV����Jκ�eW��ٝ�R��õ荊K,VNI����7u�h;>��j��7N�\����������P��͸T�lNڷ`�rn�8�صFl� q.t����B�w��a���a�<��T�fYj0�2 X�5�rtGk	U,k���t�*G�XG�����@Βr��"�{�^���3�)����b�rT��9�}m���uX��< 8�� �>��_�5��3�]��?�]�v�����2J� $���Yr��-<:��r���M�/��q2�=�����zI��	���1B
�^��lnĺd8��*�3U�X�@d��sH�� �k͙�P�
�U@���
�T?�W�$L�"����h�ܰ���չP��폛g�}�H��O�ίAq2H�u���S,�s������X��0�'}�M��T�r=�H��h����d�dZ���<���$�3N\L����Zy��b�n���Rs�!S�q���0ĭ̕�+pF�S�x�/�q����\EF�p�3���+���X@ �B���)���x��߀qNfDC���n0����ћW��	ҹ��W�!(x�����!�b�Ĺ[��\ˌ�z0f����UeMS,d	D&X6�EXZ�<��G���k���֧ ��Zj��D��2��7}�݃�ȡ�٥��S���3���8*۸I��8��W���~홗���:���Z������������<lx�T����P�a&��Q�dMd�q�
�s�C��Oi��P:@D4��v��[TZ��՝���'鄰Dd���u���%��$h�ȒL�j;�J�Üu�{3ڏqR*1k���?��:�"cS�Q�h��bYQ&�=B��Z_�;�U_*��p0��99�P���/b�8�) `�r���-	����;Shb*��P�Q�����[g�r�!�{��c�q��w:5���s��g$��� ������ �����mg�����Hl�Rt<��N�׈qW>b�V���
ޛt�<V�w~�2�����f��j�zT�G�7�?�o��Ec�6���iN�ե��-0-�C��[RD>�����[&2my��7�`���
���>c�d䗑y��U��G��	¿J�(�]D�-����v�{Rk������UC������Bݣ�nG���W�:���Q.Y�����\���9 �U����0L�H�.�L���W�Q�����}:��2�f��aB@c�Yx7XS�>[<��A�%�zss��5��ᮯ�����$�����v���#+_k�_�~=J�����8@��5|�1j�����t��p���k�'k(V#t6R?���Z��\|���x��{�fP�oFc) P�d������pԚ�cu�e�szu]�}P� �om�ȝ�LY�p�4P�E�Q��v�h���R\�{��Im���"�z:=��X񪹰EaVRG�oL׳�|����v��i���T;R� �#G�L�ҹ��w���a��~� ���y��p+��"7-$3pt�MG3o疡r���t��ԙ��?n5?�|�?L�J��������3L~y��S����w��i�|�l!j9�k��r+@/KE
�$q��)�Rry�)3T�g�`�'���[�W����suؒ��5Q������ż13�i��K�*�Y���3�D�A�Xkf���y�����b!S�daj���^���¨��Ć;G�a|��6��C�C��#N�J��Cq���U�@��en�7�P��m�q��'U�+���n@&$�z���[�ګ
R�؞$H��l������\�ZF١�M�y��0��4��\X��1����'u`��-�9Yh�_��|���$�t�[���$G�C��q�@��>�=�}f��zk�&N-����D�E\�8bp��t���V�t8�C����ƺ�ؤ+��HI�O�$8FP'�mJ��QN�3��1O�Ȗ�r��z����j��[��8�ϖ|�Y�c���LA�"&�94"�@`�-����Wf�l]V���1�@\���\}Ӓ��&��1,��+c��U�\�������b_���j�����/�y3���o.�����pe����S�z��1`��A���-�V8͞�t���H�O�M:�6�#�a#��g\��\�z�z���������7�tp���e��4�K�=`�}uF�F���1z?�2�2y�J����1��v�GT{��VWlC�E��ϐRuj?؄-�5�����s,�qq�1����b$��;�:����UGu#��N��fD�)t�d�F��m�Xq��M{~f�Ge�â��<�e8�ҹip���\s�~+DP�`�ާp�7�ے'����V�uW�^�en���I���������ί��*jvf���.�.���́Vz�OoQ����l�wH���mP�Q�8Zq�pvP?��D��3�p��]�Н��q��e��f��mb�ė]�ꐞ�B��!���A��Xe��`D�=)/Z���e�������Py���w�	�O;����F�/(�q�ӄP��B0�>�y���5N�r�&g���^G�D}ɴ��'�=4��/M�k�qFc��9�L�ܩ�D=�tA�;I�ޠ����)�A'��!���P��&f�+p��X���L����h����I3�E˄DV�R/19w��k��.���Ӏ�}�(��9u�#Y����q�cg6�f�d�;� ���YahlΙC�0��M�u��[;.�
�v?��_���\v����|՝0��Tc6�+�3��Wп�����_x����5�~Nn����[`]ղ>|�T���P+�9֋蘒���Vf��_�Q��4��UR~��T����A�����pf��ߠ[m���J�;�e]�idŚ��K� �"fAa%ˌ���p'����q|V��xh��Ј�I��01�/˯ݟ���� �� ̃�{e��}��c��R:ך��7m��Ygh�d�|5������|R�d������{�$����_%C��u��%�/2���?�U2�Ʋ�U�x�g����!xr����m��pc�0��=�ʄ[�6Qi���'v_��={��Ⱦ����5X�t��4W;��>vI��B`��ڊ�������Ui�ڠ;,���6vE���c�B���`hx'��۬斓�����t'���e��jIr����)ɷ�yY�R��ݬ^�:��n�
�ÑM��o6<�C��s`��'`��\ٚ5� &X�q�_�iZSZ��`��hL�'��,LP�'0I�R�iU�mQ��wM|,T�39({<Fy�L�^xg&���bd M:_w�K����UZ>�}'�j5Aw���{3(QxVԯwa���*Nu�vO�����0^6qw�'���p;.�����4r�o3��lv]��#g�I���cpe�+��V_�"�sՊ��l��k��T��[/N�Q���]��"�I�J�a���sQMO�&?�NM��M!X�y*O�8�z2�J�$q�~fD�GS1S(�S5,�sƯQ	�ڮ�J1�,L���I���Y�y�u]a��`��P�U����:�@ár�}Tzr��avf�� O|���<@�q{�q>�7T��wp~�ر��9G�C�m�O���z-��7���C��j}5?ǰέm�Ҕ�����#�xWrT��y�P���\(̌��1�U��b;�%�jk��hH���J��b�=��j�aD���M�X#����U���{)�dn���'W�3�t�]��-�r*G�]f�&�J�Q�k�NY|��qAM�'��gAu����@/�^���P��4���R�Ι�/׋H���Ť#�lwj�D-�"	��z-�w¬^��͓E�v!7����L�®̰����uS-�]O��§T�΢�p��s̒0F.`��)k��G~�_R5�"������a���C!��t�:�ɏy�9h؍;���ױ���fB&�~�,����ۢ'$Y�a#��>�q̟��)&ݕ;C55�eXz[GՃv�X!+��5N��1�2��RQiB���ʝ�ٗ�b�fg�R d����I����-1�ѻly�/G�!������a�	����n(k��`
I4������cMm��59xT
�;6
�����Km�D��,ì%���	"jrMn��x��[ye����N$���٢[�s��u�{|�м��vb~�3g)~K��Xyn�����_6�\UA �¬�����˙���2 W��u*���m�}g$�NI;�W�+���l$�K-�A}�/�1����p�=:'*R���Z^��������=��y[��X(��r�13����\V���-�6��&΃$׳�dU���0��r;3
�C��Q�{���g�tq񪂌j\������wz.М|��w
�.�>���&%���G��]$�|O�?�x0M���Ӈڽc*V���X�"EW��H��G��ʑ�jQ��d���z����ia`�����JY���io���YN .�%��0հ�"ϧ��65���B�)�d��������).��}��3���jh`\�G��f��M��%=���0u�U�?����ȐJ&ʼ0s�\z^�����b;e�3��@��4o�>�k�3�~r�ں��W�f_���@f������Pc�lT��}�X9@M��M�:j�T'�i���=\��%A�QR��k0�L��\��벮�R��z�F�n �
w���p��!�U/:�˕��e؁v���`dn�;ܺƹ�ON	#9�Q��3.}c|+ΪeQt��R�P�T"���8�8��I�I����?�v�:�Y��g[�yEt��?�F��V�������Z��J�EC��K��8�����$j�bYY�&S���C�#|��M`�Ɨ�b%._���v�T�
��;�?V�ҍQ��wZ��{�����&�RIi���<��R�שC5e\=o�ӻ�#�+%��&���YM��� |h�@��,��`Wh���YB~.��eW�������i��
[�jE6.EM��K�pq�s_�V�R�����Ȯ�ZEw�ckj��O7��� sƔ�\r��W0*�D�K1��HJ�F�$W��ɮ���)�2-�@"ʥ�S��E&sW�j߽],��ɹRj�S��5���	������zv�?�sCR3Ǿ��8�;�ѥ(�1�rv��������(�PJd?����4��32�r���߃�Fթ �9������*�Xǣ%V��tV ��	H����HR�Jw��!�ʕ��X@.�_Z�N�}�	�C��(zZ���r�7`��	$�R-so3��Ȗ�D|���jb��(Űv�/u��b���1���d�t^Îjً�:�裁�1������őx?."Nm��ף:"�f�(b��hYi��\	��4�@�7TC�kr�����P�E+�}b����Z��AU^5G���B� ��G��A��� ���9��� �㪎OU��ͣ^a�'mP'��WL�ɝ���D�! �)�����5 ��_-bp���rm�b��:��G��Y����Z�f1�)�n�a��|��CW�#"5'�SGΰY_d����]��u�)��6��JE���qy��G=�q���w��L�k]����7��hW�N�!r�9�l��r�
�q9�?F��y��c�X�W �����/�����.�U��)R�l^X�w-����M�rAg�7g�����|._��g�A���h��.��X^W�knfkĭ�5�
�E��]���fl�cp}f�r�ۜ�)C�*A��G���:;��w��'ܕ�R9_&Ց�d����G;��Ab�t�U�+&h'�p5����rL���Ovwiч02W ��.�E�P@S@��-��
i�z�@b;�~���Q���	<2�
�<�r�Ĳ�S轇����F)��Q;��&������#����FC1P�s�:�'K{����[�8H��E���MB�4c�;��m6��9�~�Gy-�5��2w(������.�H2�.�^��;��B�&��5���5�=k�N�����@����+D=K�}/�X������1� ��G:�<�zR�+d��~�6�zc�eP�����A��P\�i���A�jK鐓�������!� |�����#HQ��VD���� ���E�A�q<V�I�z�N,ME��(��pxK$������<��g����I���A�8 ���8���)�p�Au���%���q���q�{�ni�Xko޷/�;O�A� b�3�(f�]�+�������8B�J3��Q_�����K��M�6{�iŅ�6�Pc���J������7TC%)�W��/�6O�B>�)(�hd�\����'?\�Pq	�\5��J�L��aW��Z��Qm��B�Jfa0dމ���!{�>���ύ�.M�Bp^�1�h+o���nP�d�@AB<}��b�88?��C��fө��fG.�Kl߰Z�$���!����"<\Ӧ}�]������w�f�~�j�`2�r}r`�)@>1��h�'�P��f��3":��4qǣ�2U�_c��K��!`/DE�ʟ�	��J:y�X0�)_Ԭ̕�T䔯w!zD7�J~���%~��#?p����4���?cl/�Ǯ����(����� O��UJ��f�2�\����s���*��^�2��CS%�U�J>q�e�1�0�X�?�+�M�6�q�d+�(w21vG}�e��d�-cC_j���ZR�	�a��.vC��a ���@�k(.��9D��Q[����:�
��u�,	�`�����9�߹�Ψi�5|	>��W),RU���(����a*�N7�P�V���0�7-k��@��	����}���`�s�z�.�M�n.`��1��0����!�o9����:A�Ws����%T�D��E�_%]4g���=�bz?�p]ŋY��Z9�:�i���Z�,��ѺGE��K+�62���F�u��q�m���:
Q�"�v�>l���=�?���Ϻ]��Q%Sӑ��g�����HF�b���l�]S4����Үu������n�����
a�>Xu�"î#g#�r��n�a� C"����D��	}�!cxgET�Ծx�v#$�`#�~IH��E>b_؀����ͮYp<"�ٖ+,G�}��hb]p���\RYBsL����Λ�y��E�V����OXB�[X�E�����`�ND�Ӽh=�:�]h�,�]�l	p��>���d�%B�]��S�jn�Ӱۭ��!!2W۸�W�]�`ڡ�ʻ��W�쫿3)��[��*)c��'[ �6-��,��{SyO��﷖�l"aO�m���~�N�6�`?L�H9� q?���	�.�	a�y��T��M�^d��~�X�S��� �l���yW)6X��	D�Ϲئ��5u�}4��dl]���R}Qn�-��BF�������ˉ�so�+&��9I)�ò �;ELM�iE�B����xbEw: ��:%������.�>F)�L �t"�*�Z�v�f�}&����<h�to��H�曟�{ٿ7���f�s�n�1�.k�D�w�;�.Vӷ7=Y��Y[�h��ܯ�T�ړ09s�FPTۧ����a<����vj��q9p��M�b��eT8��N�pD�Z���6�ֱ�\���<��U@l��߼���v���]T*<��;{���XW!���ܰH�	ӧkK��Æ��K�fk&k��'c������d��;�;.@����a� 4F34WP���C�_k�v��.��!�%ϗIs5^�}*�8���ʣ�A��n+�g���~�jwܬ ��t 0��<v�o� K4�ƒ��#d�/y,�#+��b����qK�G��1����5)���fh;z��'�|�&���Y0yt�6j�K᜝�kq	�ߣ��γƦ)�/�ӿ�!VQ;���ܹ��y�Xߦn��ڎ�]�%��9�#1"��4x<u3��-���6�T���C|�Q�U_�w`Z�V��YD�9��n1�x���'�A�i�ň����j%~3R�|C�T�#�5�Q.�m �}.���-�W��)��I�~�_��>�m�3ϘQ4h8��.@���F�q���<�[ջ�pU׼lˤ��������t��<���7Fs�m%%�6oV�ս|�4꼸X���F�wm<|m3{L���.A^&�y��˛�cwr������>e��9����'��i4M��5|d����Vԁ�[��*>�+y�<����R���cg��|��$�֩�z��>��'O0�9�����9� ps�P?} '
��G,�s=���^.Eu�ֆ��W rY<.ت����E��}����S���7O�q� ��v]�CK0\>�tW��({w/��e��'L�,6Yl!_���t2��.���F� �m��#�I��6\T��o��%LJ��.�:l���]��m�^�GÇ�����h*����@�)h���V������,��s(��Z,7�%���l��i�,��m0�v�%��E>����ф�DV�>B�/'a��t~ݤ�;�d*cl����k���ٓ��Y�I%����T������7��C�i������dc�Ӑ��ۭd�&��S�ǲ�K�"��Q���c3��2�T��;���3c$)�d�x��&-����(}�X�c����*�)2�#f�k���'���ax\�wL�����ב��%���U���#�Q<��N��|}m%@A�йGq6J�/��i_��+���7m�\8�c�(�3k�`�;�D��p�h�h����:H%��m6�����o��#?�h)�?9�^��w��Pc�+�&'��/�y6<�7Kf��&��k��Qat�����0�ԏ���s ?c��]�B�CFӋ�)h�(�W�@��(�Xi5�!�L�N�6d�8�l�;����\�n���5l�ͮ>�sA{��Qy����v�h<�e���թ{ ճ4B�rDޚs�i��Qs�IT�H�s��)��q3���3� K��Yr7�����]�6�ݚl�W�s���lx���W����\2���Q�-�n�b%~�Fڱ{�z���6���yڷ��Vs��
y7MZ�"�3�`��JN[�E��ە������$z5ay�Z�r�Zw�M�`H8Q��Q��13��z�
w�
�U�j&9�q����K0za��Am�_�`���i^~�ϡi�\(�́�&lit&-9f{�������D��q�}�rf��������*�,��QH@(W�m�8ǔ�&�)>�-��
r����@�߰4�{����|(J��,Wߠ�����4`��6�����h�'����ј�\�@�ED�1�:�y�&���ez�P���_�^g����<)�)���
�qbK��jK���?����w4�<,���6޺1�?�P���P��ҙü��;s������J��P����0�Uh
��`��������F�c���wFÁ���5*��(���7v��z�n��7$�$љ���Q3E��z���4p��UW1-�2�J<�غ�|��i��b�p�}�.��<�c����R����	�\D��#,v���KϋӸGT��U6,$���6�x�8�KQvMle[��	�i�v@��6�hVe�O�I�0E[�H^���p�1\$gF��=��>�tԶ�^���1Zt{R�Je�ؐA,	��4t�G��% :Č�w�e�'��눠�a�K�jS�{�f2?ŮW�(�\�V?ʧB�t^ŭ���7W���@h��7���Q�4r&1�Y.��	��bn��We�R;�W�� ��R����I��`�qү���U5��:��R���U ��*|�#��/|�0|��UK���%�
ġ?���7����5�a�4w��Q����;=�� �H�g�e��� ��WHT
��7O`���V"�@�_.!�gS������h�宥j����7+t܊$��߳�=!� ��t���a���و�p� g���^�S�)2�JE�'�4�6$1;����:;����zڷ:�������;�B��O�g��݊��	�4���k�- ��06Ր��QE�,�nZ�i�5)
C���Vc�b&�ka�6v�b�!�MS�[RTß����:4H�4IW�]�� ,���m�}b��f�T�TV����{(HPkGóᨣ�2XA��mJ��M��n�G�����.=G�� ��J�K��{sGZ��Ơ<��(cӑ�"�$�:��&A�t�"��j���5�è�d���W䌫�	D�6;|�Ē��]Չ�P�����+�!O)�4�F߆ڞ�B-���C�@���� [��m�&j7	2�����	�lTϊ\!�4��y��F<� ��Kt��r�(��ɷ<M^�I9|t��ZLi�xj�w���,�i�8�`��t����{``1�x�I�������.�������6��ӥ�ĵ��7�1��hl0��@�(���>��Y,��8�L/19�ø����_I�Zv
5ඕq�t�GѓP��Ul2�N.X���W�#+�iW���/�����Τ(�`9��Q;	�`���0�uO�nD2Z;1��A�D�bK�A����D�n��]�Z>���p�k6���/M�.�@��^�o�`��G�#-(	@�����:�t��/޳���}TJ�Bx�pZ~��E�oa��#ͯǚ��2�X���Q�\%z!���F�����0�L��܅��Y����[�&1{�\�t�y�)��t��Jh�{I#����ò�A#i�΋��8�U�W|&�ŭ��`��ߏ-�$jX���w��\�io�{�7���	cb4�Y^�������x[WE����D(>-�5tG�]D�������%/����w�<�4ō���(<=����^�K�'C����p�0N՛2���rD.�#P�,#��6��Q��$-XW1��E\P���ŉ Ap�$�����x�>�k��9x�8�=�]�m�}Z]ӗ��S�?�\�7uJ����G�%�MU���g�?بcHS-v��E�J��V��ǡ�u�zcCr:�2���\N���h�m���ԙӓ�֡4�_�#��:�r!�p����u%�3FG����zcT�>��A:�S�e]����YR�-!Sx_��Rkj"�(���i8s+����T
�ݴ՘���$	����B��;�����ct!+��]5>�؞s/_�b��A\�(���D/��)��0&A��:8F��C���6�f{���n�z�TyNi��c��m�~[�<��aQ]�� [�(Nu���d�bsR�����q�]�	k�1�g������(��E�p�H��<�ړ�*�)�2%����,�� 7��@�|D~�8V���	��_����~% F/�~�#���,M�:g���!A��"+�7���hJ��S��iX-��r��Mo;	��&��U�Y�x�ˬ*C��)AUC��f(�}�ir�ce\�H�c��OHC��7LRo��@{x!�D@���dӊz�8(�@���/��l�qw��7u��Z怃����}2�%Ү��j�k�fWj\L���t�D�||�a͂px��t�C`U~J��/�8$�I�w��/��ɷ4Ք�������2�%.���w�F�~�	��h333P�lw��#z�J��ơA��Jc�+?��ݰOYL3*�< �˨1��#��"i���!CC�!2 �%�3��R��|���ԝ/k4��T�z�����R�{�W�6�������9���TO�c���%]l(��lhh���;��i��r���1�+�
���5zC���� �:>��5�C�vt.k��R���k�W�7�A��o���'��2y@�%��K1B� 틿�!����;³W~VE%4a�F��׳�Pu-���Ԋ�4Β}��LO� Fw҈Y2��+#�����`7�Br�D�!�_�D��0T�} EܻvPi�i1�u�b]����,eU>�b��T�T��n>Y�4���ʇ�T3�=�W�9�YK`r-�޺�(8�z��q.J�
�,����o�D�P�K��`}U[��1��O��Q�vxt�Í��fu��[P��ڄ��R��	�ױ��I��[���lW��'v ?������f�Y�Ƶ2�Jv�V��P���,�	��e�d�Ee�m�!H�\��cO�<q��J96?�;jK���#B�ɻ�*LY���L�n�Y���(���C
B	vjiuF��S�Dk	�5jH 0�D�@6��;7$�T���e�d�7d�ۂ��.���Ơp�oF�#x�ݘ�Ǹ=��~1�!&�0�8�xPV�+,X �4��HJ��>ϲ�:�\���p�n����8�T���$���G���j���m�*gV8��9�<<����4���n�J70�D��ݎ�7���r?�`� E#�W�Gw�y\<p�>ڂ*�[�*�P�O�̭��(d�?��5��J��dcDȴDS*� ̷-�"1�� ��H;�e�z�
���h�:�c����G�<@vF\{�x��P�6��h���W� g�U�h��G
x��} @�xG�>�p�(�;$ oz ��gP�n����<�w��4��`�Y�E2Ypל���Q��D$�����ML@;ǩ�\�x�,�/���t[3T F'x�귵w&YG�LR�Ɯ��G�E�Y��x�e��m���^ʊ]�/@^�?i����/fgCQ�a�EHL�fWNe���S�f]'p �����xs�~���S��2C@�q��v�pu�K��n�%�
"��.IA=P���O�&�� ��56���e 1\k�d�4B��!��]����}��
������	%�Ig�Xe�O1�m��2����������pX���3�zgn_�T��� HD�.0M���ӊS
ӰJ�Ȓ���#��N��b��6���+�n/}9XE>�`��Z1�,Y|x�v'm9�� v���v�+��(e�ѣ��>���&iRD�	�����n3	p�� {u9��
��.�^�~�9_�EfT�{J�B0�߰Y}T�s>�W��� �7\@�7��U�p��!{�?C�^�>��#�[��~T�e�[/~9�8n��k�����[b��Xh��XJ�J�3��/̜����嘼��/�k���H��V�ü 1$3�-ɪyeXI�ZPY���:OiI(2�o��9_� <ա����=�=i�n��J'���b3o�x�0�_D�"��)� �n݃sӐ։�EZf$eߚ���	�ܚGS�r;�%1����?����]���9Q���������Ż�A�h�?���Y�r���ϳ����Ql��T'���>��,ʄt /�F�"�c�%�+R0��pƫ+��!�yd���0NO�>�dUOɦ3�n�3�)�'��1�ZTi�k���C�$�
�/����;zi8eD���G�fZ5v��9j*��?iW�Q�M1��uQ���7a������Fz��@Z�G�(.<�^�c&vˠ�B3`j����C�]ޡ����@"0��c�)�`��Yq�ZVMU�EX�A �%\��z�瀼����>c �fH�#w�3�
��ļ#��m �eh���u��],��S&U� ��/1�����k�~+V�ėB�S��T�Ŷ�3��G@C�F5�ڙ�o����=�p.�%6�V�Bu�F<?��HD���X�E��Qsx!�oGj�N���i�����N:I@�&P�6��TR��Fv1��j�m�VOG`U��ю,b�U����H�d�:ϔ�{G���������H�z��ڜt7�q�{����Y9��)v��*�`�{ԣ�J �G��;��/�z�,���,�,7�e]kkF)��!�>�fr���on�F4م�~$�U����ɓ;���67G�CGx^@A|���K�� �����(۸L�R�zEZ>p��@����|_�	�ze�и�eM_*��K\?/�-�G֛֕4m1xW�~aK	��M0�F�-3����åE��='�%©�����>{�ߵ��^c�һl۵3��wɝ�����/3sD|T�p�����Z'��staO�)����'	���?B���K�HB�O�U~�>��v-��gon��_���
�}�O����ֲ߄N'���\$�>��0ߖ���>f�7B="�O[��k��r��<ˌt���[v����^����[
��'#/���:ְL�~6Y\�	�>��. �c�세,E���ऋ�4�:��r�����z,)�����A���r�z
�# `�t��Sۻ�ĝ�;i�?LsD��P�x�a����1�lN47uNePx�s�l��+���Y��
M��ɗv���G=3���0]ٯiNt��	c�.���}`U��"#�>��ߙM�!Z
U|LT����\��* �nf��@ť�A �Un5t��k�s���PA�_��2�;⩂���y��d��|��Q��`���lx��h<˲jihl���Z��v �s�ފp��n|�/��s����Mǯ>�\�q�9�8vZL��B��� τ�C)i�5kσ�j��v_��ض�Z��4bϸ�EV[�[���G*yq̺a�"n����L�:��̀/���}��6�� 欦y�?*lrAWY<m����_T�l<���U#Dr,/�6r8QY�C}p��2�jOfF3�\����-E�����Tb�7�ʹ��ʉbj�R#x�08�W�V��Q]�f��������{QH�:f��1�P��I�?�j�U<�h�l���~���+��Գ:�������Y�Zgߠb�5�[�^@W�\���²������e��a�5�,GDI:&ߡ�"�l�>��L6i�aoM�Q��I,� ~H#���ښhҲ�j�Ց�U������s�#��Y2۴�*~��O	ز��4�8)> Gު��̷5A�K�o�o��&��T�8q�H4�*7��_�ao�zJ��b�U�(��J��5��(u6�_��ȷ�5ٌ7L�R�
gR��_�e��d���vK�P�}�ލ�ܩ�g{�ɔQT��������7���{��[-4��X��jN�?~�BA��^�[D����;y:�EBm5��!���)xm��"G����	���yrd��6����@�T/�q3_��Om���w��>��3���.�x�ĭ�fȮ�,��T��c�L�9 yE�2�Ev�Y^v��5)���r����P(���[� ~?ag��>�R�W}�J�����1� g���Fy����w���B93 ���������]��_ճ��	Ƶ�
�é$�����ޛ.�n�A�J�	6`G�3֦�c������V�u�L�kZR�\>%��$-�&��}����EȣS�4���*�A���Jf�N�>j�|�%"�>u����ԙ�}�cp�NV,��_���h���;i�
�!�sѯ����	G���-��C��v���s�Q8��7�;�X �U�~��s����w���c�����X
$���kRK*��W�s��@B�|���))��ėPn���qH�!�Q���6-̧�'Zo��:����9O+��'�w����0��'�h����pa�K�����<����U��fW���۹��g=�/�t5\��9d4��g _�f���A���o=��K�f�8�ȝ�=�[��@Рe��>�hG����K��+�fU���FDM5�dy�My�ub�ݹ�Gf�o\��*дgOݱ�D��r�� ��3�!
���b�-WmF���>|g��Fǘpd�zm��q'ك��[T��j��5^�-��������D7�~���c�}�TF��H���b����!C%�t����
���S��뷦��V?b�n��1��;n�=h4���R�FoęSP¦�U�9&k}zկ�l�.@�Շ���ƧX%��Ի�}�.�n'�dC4	��B�=���-���[�U��zhh���Ɨ�Uh�o`h�:ō�!m���M�yu���hܫ�L�}V ��-�Mhz�9�T5����P�5���P�xWHf]
a� ���Ճ6��>2K�\\�'_Q����@�vy�HC�R\����4�
e�X��ɮ�I�8��a(x�Wo�ɸ���>b6AyH3v���A�xi��
IFSFˤ�J���SU���)����pvL�D���"fd�X����?Y�����}��5�ߺ�;1�,¬"-��5>R��+�����8ؗ�����W��M���L�E��� Jc�
,M ��r����o��>�N��W3=�5,Z�'NT�6���M|�F�N@b��:i�}o��ѡ`'�	����j������	m�Cy��t���o��>��MvV�n&P�M��=�<"rm�tKQb�����8�����d�)U�c�2���X��8����f���W������qLBPU��	��r��"��\�O��d<Y]m�̆Zc� w�h���OTh%����Ռ�E����ɨF481��[�p�(D�ׄ:_P�e�rK�;�=��0���B��r�s2*���3�����!��bh�|��5L��s{�3-���թj�<x3:���-�R����Ea&������eB�+�c����>�T��7�C�Kk�wi���t��)��%�~ډp��3ꆣV{z+��Gӵ�O�̵)�w��fft*\T v��% �ҕ���8qt[���Tsgc���K�?$��i��Z<6���$sW�@�x�|�c�e�sR�ޚ��a2��#Z�go�ep�!����,�$,FK��q}/��{��1�Yb��h�q�Y���u��BY�Ԍ|�'!�Xz�8}���K�lv�nV��B~u֞@H�c��Q���+n�陧k>x}5<5�+��t��N���Ge���b[�M�Y�����ޅ9fv��!/>-7�0��J�yz��=� ��B�9*Y��j�Ku���� ���9F�{��ӰXgǽ����K9ħ37�|p����-�>�I<m^Y=`����(8}��޷;��rH5s㍀5�x�p���4+�y kjf�0���p����l��r�3��x���_�
��}�@FM�5�~Yg ů��0�b���yv�7I`�s���h�dou�8*���f�����V����]di�n��Ђ�v?�;}��*�<����ùE�e�R���[&'���X��#tK��.�T�Cc^U�F��8)�F����nM��,al$3��_n���~�G�ͫ�9�x��'�8p�q����s򳑌)��8�J �5%~:��Q�Evs�C�<n�fG��gsP}fZ�)�V;)D�i���N�扏u�p]�����DFK3�
|+Hκ�J� o�eB����
2�g����j:ڼ��@�e�e[3�<4N�D*њ��r�s�*��}ɫ��q`+c!Mp� ��;�5U5=�Am@�Y�'�'|*���֍�x���s �4e��E�}��1Ho9$�ZP��EF�����0����,�b��O�d�M��d���`��h3�O�Q+�u��`�����b�+�hv�-ʋ��m�W�_״;��V��1�I~����|��+֥����K�K؉��F�0���
	��I
G�ē�����*�!&�x&�N�#?�nS��_����K����`#�Ǐ��k+I;,������jEj@	6^m���cw!�w(�� lwK��i��&OM�D8�D�@T���a\�ݚ�F9P͢�ל�y�\��k��`K�٩�[g�#�E<e2������GЮ�jG�W!��淚߈�Y�0_�A=��n1UJ�o~������y:-ҕ}�R���O����2���a��8�d;��^����Z�,��䅯����_�Ӛ�+��,׳L���<x���ʘ
#�C�'�+�U΁�BJH�_�Q�-���[4^B�;zs�ł�m��4f�����|�`i��'F����x�[HA�U�o:�vOxz)��V޼�eA:�D�I8����b�����b@A�5H�g��.�Gq��wSu��[��%-e� *�
�$�U `?9��7y��r��ŕ_�&�1�.��^���!�@V\35.�ĄvV���4N�^r9���
�{H�� �k[�YH?>C��l.w�&ٌ�5�i��%���C�������u�"���rT���C>
�����|Q����`�d�l!��q���!�IE���|�u�pjK�?��~$�aC�Dw� vC���壓��!�6p��Q���)^I�V*�{����7��g��������ue#m:rEr�t7��H�.�Gq�%�#ߟ� &�vmI�O�)�T�v������H�`��N��>�M�!����7��nL��>v���3*P�,�wD�٩P��W+�B���[���/u����1���[�F�-��-Ĝ7����6�7���P3��m��8Wo��]��m�!H��|�aj���?���3�b0��Y�Ľlu,�5��ʽ-@u�P�E��O�����c~��W|��E࢚�u;Y�F���!��A��7&��8�������_k�b\*����kY	��������v?w�����g�c���f0����'�d�O���S��Kc"Y�>���9N[p��μ��c�.�
�Z�[�F�f,cF��w�u1�R����o�����i�Y(��y�gq�ϝ��q��]1 �16�M-.��6ߚ�_�"/-\#Tm�[�����~Š�����Hz��\H��+aQ'��;!w߻oлE���Ă��KQ��g@)�_Ζ�@��s& �벛�C�|�J����d��!�z�!�)�/u�[c�`W��k�"��+D�"���v���ً�R�]ΑtJ��!���f8��3�q�#�8c�����yFy�~Qs��tm@���&��x�)"�	�<��q�iU�A���=nn�}���S|������<r�K�[���<)��?;i�yRHx n�n��3�Ĥ��j2/�>�)|���}�k®��B���k�H}w�G�,S�>��?���þߥ*�U����c=յ�I~��OGP`�@ȧ_|�̚���)c��Ĉy�s�){F-ܚɡj+v���<� Xz��T��
+�C�����I�R7$0h:�S��ю�����;j���G0��_61�%|[ҏ�!)5 ��:[������s]�4>?N`2q���Y堁UgQ! ?|!�rƪ��
��H��5ׂ�hN�j�ݏ��F�����?��`v��z���3�<���6�fg����neCu��A�%Vlf{ǩ"� �d/D^	m�������p�������m]�-
ӽЂ�c���z;{������cö��<%d�fZ����uy�ݓܔؒr��Q+�w����R,�	r6+����	�V��߼����*e�cJ��2��f�N���d�� U������ENY^�J�0���adev��h�ϭ���D�Q�ώ����ZrD���dNuH҉��$�"��M}P�P�;�a&�2�3w��8m������{�+x	<M
�8�*(���'x���U-\q�-�%�_BJ(͝?o1�b�Y.	�6���0; &�,�2j���
f_��.F`e�O��aבw�e��_���O_�p�
���r���X�|p��aaz���pbZˌ�}�;2*�9�q"������� ��8�)�#je��"!�H� �Qz-,<pL��Xfnගf�� �)�D<�F��d�����O��?t��8@s�����@e�n�"k���3a��j���0�4���MZ��2Q')HXғ=]�1����"���qC��Oay��rf]
G���_���<��c��pU���N�eڮ$�� �d//{�^��xؔ�N��`�Vݖ�>Z!�pLap���GZ׻��j������G)��=VD4-u� N�@��d��Hu� K*TB"e5�R�d�r��:Br�����cڒ���:�,n�D�U�!�Dsuމ�s3��q�����>��w=�9'�?��o���Wve�?�l<���̽�x;�hR\y�W���N&���tyC��	���@�M9�����yr����v����C�����
5i`1��^K�i/5nN�{���AF�� �,�:�&��"��z�8F��G�z �]��ʿ&inQ��	���z�y���+d�@�T��K_�p�i�����|�B�����$� �*D<��xi��1A�Y�^�ȝ)2�x���F�T��Z�Y[���OͤA��Hލ�nF�4<Q��������XT�//�:�V�Xə,�� �DWt7^ ����`��ڋ�f_K�q�t�^�Sʟۚr����1k,�B����� �(�nW-x=��[�!$`/��Ou�L�]�O��T�g-�>u���S�|����;J M�m8��XO2��2ei[�W�"�)�	�{qm,�G�S��ڶX<��
4��g�W�#�R#����c�n�C�s�`(	��>0��`�l{�to�|_^�w�`���T@On9b�N��o��z~Jyl��RS�����Zv��bX��%l���}̒��)���9w'�V��{�W��F��0s�%�"���:�L�o�q�ݐ���@�3�

	ي������c'U�����JQ^&�7z��k�ũ��̕�]D"C���Q��Q�`�3c���:�â
,�$p���ryW�e�NǏ���n6�OM0d�����Rt�H	�~�ڀ�"�j?������"_!��zL�@.�����!+]G�g���rhs1`�\��%Cu����9�h����笱 zp9��`l�#����>�F`yPøF.׉����佘�p��\lꗤ�|���T�e`�,>}����0-�(;-���"{���Rɧ��L�8=�*��0	����A������1�yz9L��}�)�Ϝ@�/��g%��@5S�9���|̌��Fm�R�;y�j/f�-fC����ýv�F�">s��
{ٜ��`��6
5�g��t�Fڭ��G�Y���넭v�_{l�V�i�ޯ����c���&�A=��[���鬠�����y�'�T�@�e����G�~a�%jH;dr *r]G�̃��	�{�^Nw�S|���6�� cv<�0֤�9�Pm��$��5����ږw�s�nu�V!pg"+�r�1��dv��4�f�W2������h!c+Cg�{1a�bA��">
�*��o��(�Q��S`V�w���yC����R�����C�d�6��CN�4DR�[ʕ��o�}��}t����k��|<sv%t����_"̐���n!�Nڥ;��P�k���D��mlֺm���*uZ���9u�s�`]� E)���^��h� '쭉\|��*�&��a�$�>.VMdK��t�x�k:�V:t�DX<�s�i���p���v��!c��,�e��!2�:v�����|/�m��g��Őhor{0깾h⢥�8�f�j��i܈���{�m��%"a�6
nF����^P/�MA��촓Qwo�5�\�3��R�	@� ��2g{�i'�H�ŗ���P���a�^�_�w|�Kǆ�V�{�g�r9��]��|��;A���5"�+rA��7f��R޽�*�,�1|��1��Y��SM'ɟ�'$n��b�٠�(�qH����~9�=���.�4��`���,j��UUT*{#ty��I��6;�W-}��Jȏ�G�N��o54�M�K�����V�m�Z�0���첌�F,���=Oc�m�����T�� �YN�Y��`��89�7�.-΍_��ѡ��k%�:o����ܷPjO_R+{��_1n˟���'�����@�O(	W�FndS)i*�3�1����2�3���L�ȟ��K%�Y�!=��&�Q`��o.��v5���ٙ9ʂ��vCJ�[��w���#��aƼ�	
���ȁ8M6�ÁWƀ���x�i5�9�.E*�!�^y�����V/��j����Vg~��TA�'�3,ʶ�C�D��|�>iq`�}x���n��i�y����j�C��0���Y_��h�u¹�I�`�FK�6��5�����uޢ��g�"����P�ond�����Z�MrC�gVђ�ꗊE�x��a9D��V9V��Nl��W�[褁t�o��7�ANT�el�}���8:����X�9o���s��	O'-��h-�%���|����3�E$�"U�_��zm�|i��`��,��vkx�d��g�v:d��-�w��R� _�V:�"¡��H�0�Tb�u�W�k�*��H��oe5�k�j��F|�t��B�0��E!�����AA8�	{r�
ⲇ�Їgl��G��f�T�oB��8��Ά{@$bA#c�6�j%l����7��@����*V���䣖�����R�vuǛ���s��x��H����C��}�]�!9_��9����agt"-=��t���$� B�H��d�Fq\C���l�Q /357��A%Yg@R����R�����U�������hwo㉮W�e��z鳈���J���fpTJf��)��7S�����$矽���[�V�֑|��YԨz���c1nXO�X	e�5Qc]?[�eu; ��C�e�#�����֗�FwOX��a��G�g_C�#B�bZ���i�^�J���S�!:R?�	>�"d�[��w��E�K���ȓuꪥ�H@�z:�73od M56d���e�V1����CX\�0�L|j9���������3���lY.Z3��n�C��Ǌ}�-��^��'Z��8'{��H.>�m�����{���>���@}2� я��#��K������>�mmG�
N��s�ƈ��[��y?V_Gq��;��0��V��b���Z�Q@g�b�R�c$�Mv����0I���`gޗ�8����[KCq���)�`�w���&�x���#*;�t,�7���Bt8{�{�$Y�aC���؄�c�ѬB#���a��KAb��Z�.�O��v����J�t����<{���P�Z��Y�i]d��t�oS�t������)Uj�R寧r9�Xp	�;l�/���i)���e7g�޿&�vu8�\1��X�xӮC�nx���ƻ��9_�p��jJ�!���	сR���.����|�� �W�x�Y���Td�kXmv�ο�G
Yy�
�f	8y���1dT�u��k�v���Y<A(��Bo�������bq\�A�H&-�h�J0�&�ʲ©��!����⊤�Z�jK>l0�Յ��>9}Ab5�*�)�7}�������Q�G@��-.�r����rs���^'� Gї�SC�r{h��V�E�����,��x�n]�β��tUm�m����"k��1�"ӨK��ԏo7��,�QO�f~�c��1SZ1��FWm:QG)�"�ڬ�E�hY���	g� �G���p�ƏzN\��NGj3N@
�B�]`1�Y]���f����>��w����dsR�<�2�6�����Y/�aˬ���N�ԍ��-f�X�Т&�fŎvp
2�wG�q��+q���
 Ύ�|t��ҳ �Q���/d��H�aaI.tz��fZI�R��e�"��D0sF#9�e��]�y]���q��PD:&���|�3RR��S7H��*�~7'�V�	�{��0�Nv���Xd(�����,˄:��j;5���Ȑ�xI���9�hu��,�bO#H�$��B�z���a�|M&g�c>�RЏ՗��n��^��:c�v�aN��Ә�n���Eih����sd�r�)�Z�䴗��/��M*��C�.�E2<d�ĥ	�@,�H���{R�@�̦�O$�ܼ8�NT�\(ƺ5DYnHFW��V�2�{dދ)S��K?_㤝T�ʱ ���e���������p�<-�����@Vѳ�fZ��؟���K%��Y�n{�Zl^�o��[��Ԫ`i�#D��Ed��E�x��L�[�[���~�9#甄���Ws<�%�C� "U�=������2�ެ�Ox`54������%��.{�B[�݂:��M�2�?	��J�;�O��3�}�M�J�ST�=C
:!>ʁ|酗/
¯B��q�6ѝ!�|����~�����`��+Pض�Ӕb�%����~G�
惃ps�yQ1d�#6�~�2�Et#��3e�噠QӾ��';�R��~�ohd��[��2����Bb��?��>���N{���=��^��ߥT�mS/���,2`��Aw9ו�g�3S6�L���;YO.ί�����1#Ű���T�MB�z��O~�\4��<]�T�I0~"�p����_9�?� ��k�Ue�`���́�հ�1`ب�7���fj�x�!�� ����㳧��\���w��מ�D�¥jU�T_Tg�7Z���s^gF�
�0�ׅ\���qg�zi�E�����+Q�,�헰���/F�ަ�;]���C���UI��ۆV��t�'MIdhҹ*����2��|"ԃ��\$��a���T�eKr�ƚhP����?5ªl}2��A:���6e���"!�I����$�a/��r&��^����䑂Qf���?�cІ��ʙQ���&Ag�$4!@���}%��0��#:�l��bj�n�RG윐l��e�z�0p�{���`N?�23§a���D� T��Ŋ9�J�A�U�Z4�Z�Q����{>0�%�Q��/���Z@�c�J,����vz�����{�@9��k��I]$O-�����,�/�ۄt'µԺ�s��B���t���=q}��a#�J7f��J���`�3C4��T���(oJJ�K�y�!���Eh��@��;��b���k�te"���j�	����K�D�Z�?�'�����z�'	�Q�?�1��R��}A�����w��6�0������k��|��_��I��߯|��Ͽ����,x4��i�9Tr�U�G5����`" }�De�UP��j�e�>DBj�1���O���OL���-_�-�{��E� 
}I�v��I<���\�s��&i7i�^�&p�0�ָSC�,Cg�o,{�\Y+��:�v���P�}G��8�	��P�)���`�z�A3�U�=S�&F�4��j�*�+�Z�ױ ��F�л7�ZS�W�V9pm�Zٶ��CW~���X�uv�ZQ)O2����Y��`����Ћ���	����G���G��Br�û� d꫌�ϊ*l�?��9��;X��O�'Eo�{#���9(@`0��S��1�k},�d��Vb5��?��=�� �S��j�o�ZC5�V����j/�����B�����+g�}Ǉ#�?�y�x�0�vq�/`fֳ��k�C'�N�5v�5nrs��~�G�d7���"@�j���m&2vo���t�M�3�qx�`�dn�P��,��uU��Ve퓎;v�ڈ���������HOk�$��p�{e:ʀq�!,L�->;�tѰ�v'I25�;��o�Go�����뺼��}$ȇ���@��9�r����Ӟ-_��t+̍o|�0X������n,�d��u��D��?{"�r�ܥ���b��V������,av��PS��+�3R��9��fS��4Y{e/\��%��~��PJ�
 �Q5F
�Ttї� ��ZK�87�q|�FY�����'� ��<����u��<G"!�j>k�(�d�v��7W �AS��3�q�N3��y�o_ܩ=�L\��\NZ�+�Ӕk�ht?7˕O�w�ʪVV��}��&��`��QYo�Q���w�C{�������{��av�]��_�t��Ϭw-�&<��}'*JDK.���+2��Ț<��5ʏT� �����8ЋD�3��Taj����c+�9ݟx�'00���s��V[��nY�ZE�G�xAۏ�Ձ�i']��ha�HO���/ɴ4r�w8D��>���_.?��J��7�m�oV����mB�~H#��� �3%Mߑ,'��e?߰��)���OO$q^�{Yc#�h��6�5Nf}ն�� �*�=�>�s���R'Ǐ���^����ݑ	�=�G������~�L����4H��4�
��v}�
��_�m��v�����N�k|8_)U2�	��=
2HQ�Ka�z@�+AwL_��R����7�rr�_:h]#e�>��l���D��瑏(m�@��s��*�0�*yX.ܵ�� ^��h�OzM!��a:����Q���A�W��j�Δ�����4�ۈ/=ܭ4�I0C+-��ҭ�,�I��'hu)g��b5��Z�,�����?�l-}��J����0B����e�Ue�V�O[�T)��Ox��J��8D<�_HT���������ԉ�R�s=�6$��؃Pߘm6��݉q��
�-֠y��S���j#�E�L��R+U���EI~X$?����u�T����Q w��������7@�Id�����y�Bv"�������-i�]�F�Sa�m!��N�\%�EB��^[�Apڠ�!�e����3¶.����]մ���_X_0��!*��ʠ�w����9P�L��E�,�m�(�
���ݔ(b,uO��*H��Zf� S��!�{�>c\�w���5�!�Ye F��!#^�U^w**_�_HWv�&�Lܶ�9��i��l��h$L�
w� N�
��H�������S���Xy?zb����O�m)U��B��h_0}�em֒Qu��������%���,K��r��)R�a���8��|��X�5�����5����1]Б�^��g���?��>�q��'$̵�6k��O�j�w"020J&;��A>.������J9��	a��]�3 �݂s���-y�rIL���J�4��^��Q��!�,�{�)Sz����M$��粅�X_�s1ꉥ�ٮ�Wy��2ђ��$V�tU���B�Q�-a�6��C���1~��ͺk�K!P3���D������;=�V6���_N�Ee�Z�;��l,,�J���E�2~+(��B��Wa:m7��v�+3���`��Ԗ�!C0?M
�ݓ>^J���p����Z^��ApV�bE��Z��y[�0���HL��h��A�q��bM(���)�V�I�A*[t��x�C������ �%KH9p�D��[3�;��d!�*��Jcd����M���`D�ٻtG�Fg$7X��)�;�u��u�MҲl�*J��^�&�w�``)c��8ŵ1�$�e��j	w�Z�~��Zq��}+R�o��=�ek$�>��4t�y.Io|�	�����g�~y��C�w��/�	 ط���Wr%p��`}c�M��'�]R��>�a����	l~�~И�3���,�5�;�� C���B�"��v��,�F}'���0�9�����",����S��$+�3�{bF�c�`�4��k3Uj%
`�Ql�C&<P�}VEn�BZS�[&r"�H�1I�l��f��B�jϑC<$���4�]�>�3\��3U�6�O8�~Ҏ����t����J�����OT"ثڻV���9���!�[���yfSb��(xӹ��)eltE��U�b*��
׭��ȯ�T�c<�N�+f2���B6ި[6�/��I�?���`_�Oﺟ[���\�^M����A{�����2��(����a��bM�'�	~2�(�t���B������bA3rI���6���*�J`�@9���-�=��U����8	M�u�8lB�J>�f}�o������g����T�O9瞠|�#=��� hHT�	�c���4���rMW�d�
��$8G_W�2E���%���1���9�͑����H��t�O�C�J�	���͌e�bd�U|=f]�U�Jc��4;���!����'�����&���Ơu�8=)�{��L'!�G�zE磃N�� �k���z��D���ZHB���:T7;-�4�&֥m��7�q����v�~i�%�t�	��>�1&�U��!ʷ��"�fO���n�/6C�<̵X��Fq�j��}��A��]$�u�������?�sH՜~�WF��0L ���u�o�	�0��z� ���@�FEm�0������J�T����A,x {i���h!���/^���s��T^�2!�2�����@���p���l@�a�-�K'�s��l>�]o�Z���WJ����=�-ѻ��YC4Ō�?����y�fr8|�����}��"",�n���`F8F���v�� 	Iw����œ ��C$8�!3���7��4$5�ǹ�P�p~���厀l�+ّ׆k�˘;Vn}�D��|���Z�-!�J��i�#A@��dJ�ba}b�b'8W���ɮ:0"�����U�RM���!%�E��kv�=q< �gr�����5���DyĲ��wp��������L�֊����x�k�"�ȅvU�wi{����JS'9e�O\#ŸbqQ{�3�mp�e��@��H�����Q�Ihw�4��oت������&�O"�z�������g�H�*$e�-�6Kf�� O�.�t.���9���'�	���:���>!s#�d�0�=��O��d_��a�{TDn���%z��Lp���[��*������h�^e�P&�J@��#C��\Z����}Gj�m�\S� ��҆�lvFZ�m�af�M�,Gy~�L�����D!q������-#X���Έ��_�@Y�.[���x��t���jBp	��_MUJi�FA�3���^~z�MPe{��x?��~Lm��C�4�3D�Ur�ֆ�D�d��nn@槈S� �4�z�K��#�)�TP�!����R�����[�rr���Rz��Ag�`�S���I˦9�'F1��_�n"X����)�9����/�*�#i'�35iuk��c$w	������9ﳎ}ԋ~��s�L����Ve�Uf�9&���S��O�O���AU�Ě��z���K����PLe��W�H^�~�����y���Ǽx�naBj&���14���7�=�e����`�Ĥ��C�0����-�}�� �������'�Z �S6c��[o�TM�:�t�&*��%�}��RV��4`�D�t{\r�ݩP\D#뒛L�LM��\%+�\���_S���2�t<T.�����E֙���"F�Dxi�)�A���K����������-ˮ���,��3m�w���Rjn'�)m���@��OLX��]�!�A�>�^�w{���$�*�WC�v_v�h�6�j��0�WJE �?�*F���s}�6���%�g��B���[�
�,uBM߂_R���-|�U����y�20-����Hn�x��L��T6�M�!v��j��>y�ԇ�J-
�ox���]��4��C��`�,S�?{K����ZC��ی6>5�*���rU�'��QerH���	N���b���]���{"q ��e6���P?�9�-O�f�(�g������i��B�b@� Z��]�����PD_�ĩ�]���<ٞz�Z+[?'$�9#�UT���k�;�ӐS�|`{}2�d�ʀ!����Hc�Ӡ	�X�/Kx���[���&�$e�[l?^�ʿ��i�'Bݔ�ܐg^��8�[ǌ�K�AiHY���j�p\�[\RV#��3#�P'&��|��Ʉ��������h=���n��"��&��|#v*d%i�b��@�����C����={�m���R�/�]pS�q�83�&�KJI�����wQ#�?4�6��J�1������n�P�o�����+�m�
�U&�J2݋:!��k�8�ƧoW��oH쫘�}�tZ9ݴq���&�~��MW�82�O��Q^�"e�>}��K��8�w.��:�u��P_3�V9%:�����cf{�k���-^q���l���5^���6?�O�Bw�t�K#��Ƀ�[8ܺҁ����\�p\V����gH�[�C(נּb`P�8X���둺�Z�T���E���X��U)� "?٦���!�Ko*����ʌ���֛׫�Jےw���^�QB�UX�{cR���Eԥ�F���W
�7�ﹷ�F2���٪e�Gʖ�R��'��d�+;�c���&&�Y�����B�\�������v�Q�Z�LqC[�pF��-�:���� ky�}�5���J��rغ�
�-�:���y/�����?4Qew���ό�1��&�eՆ"��"�1�Wh��H�y

���X2k4�Bc�m������ﴫz�T���y�ÿQ|+B)d3���讱bpkz���D)T�E�ae��0��C r	��jK	�v�Tpd�M.Ƒ%��.�ș��o�Q<�"w��صzi:C:������̷L���Xw����t����qͨx1@�"#֬���b;Y�yJL���5�C�.� ��6�d�H��G�O׸ ���]�߫����j)�� �����0s����hFι����ꟿT�:s��3�-�#ep�;h�N���̬���	Yc?�1�BG?Ot$�kxqw�"�������!��H�$��t�}'	�\^Q��s��
	��_ ���jw<9��s�-��!W�Gܕ��D�M���A�Y��.1���&u��L@}gl~av�٪b)a1)�.��?���V#Ӭ%
}dW,֤/��O�jO�L�U7��D�#��e�:�l4�����;���}! ���}�	H`
�\�ǌ6R��2˰*=�u�sE�i��^���pƼ���	 C)�^��n�W����gw��F���J]���/K832�'e)A�o�KlPA�䶹i�=����~4�`|m:~�ʅ�ON�Bt�A��g_�Om�5\p~mp���nbpoU�#_�f�U0�k��O�j�d]�7T���5�;{M�D�Z�����(a!�������GV��@{�i��W�_ >����cuv�����[bN�^zr�pV\=R<pL�E�8�6�Ĵ�����sEǹ�ő�j�5rX�%�"��.w3:�b;/��
��6�E�p�4��Ho"�}�$�cl������lܒ:v�E�%�������^ ���SX+N\~�L���W���*�-0}3���	`?�dj�?�d��#5������F�]�/J���"䅔'c�O6b�
ӑ|[��3�j�~�%�в�\�"�J��B�-A2:e�kS��i�y��p�8������[��.�x�G:K}�+"�z��[O�N�%�������a/;��q#U�ᒅ1�Xw������in��M��O6�ݿkǤ���,a�:z�����蕎��I�r�	�!���K�Ő*�8״�����|^8�{����H�}�����V�J��=��	Z0->ù��ߴ���_>�Ȼs�����]�s�P��3���:'u�c�v 	�������@�@n T��ۙ������K`��裀W�O������S�$`h/Ո#�e� ��)?0��@�N(���Ne�a�9=�I�� �Gԁdb޽�UX���}�j�V����;�����D�����F�?�[	`lmh���5V<d�d�p�!e1A˚�,���b�,,v��gC/D��9�=�����DAb~�}'�A�0zp0h]�	*p��
5��yN��J�[�.@���i?˖a����{
)��E�ͯ����v�=hT�2	yA�`���$�S���J'�.Lp��|�&8�����\	��_T���A�a��[)0�����ˎ�=�h�(�H��bI˾�Ug��\��#�\;Ϗ8�x�t#�ǭ4�(���K��7,�"��!������hYD�h�#��]���IR��*rS����m��Y_��ưr����U6񘎀��f2�v��W�?��x�˽o-�Ȁ8	"�q��~�A%�iH}Q�H�,no�g�IHH�v8V^Ԍ��� M}���}#��~�<��h�KmW�K84S<:�V

�UiM\G�0aI!�䓗�ݰ�x]��q����VJ#�B1�^��\�c���`���r�����E������4��{�d��V�kb2P�7z�Y�����-PC3��t�WI�D?��X?����0x}��*m�z��Iw�x�S7�\��i�+��hL�Ϡ��ŚV|G>�D%6v���5�qU��k��of�ǡl�xO���% bt���c�.��ő!�@vm��q,��)*W�U�j5{�y^m�6`�}��֧�__�יz@~�羺�,Oi�%�����,���jk���FD�k�Ǯ�e�@��4��VΨ�o�Mhw*�oM=7�>� 6*0�iIb�;R���kC&���CQ��������`��i�4��0$ 5�l�
�����6��ή�<�&L���C�-��J�^�Q���6�(���f�*�N�nS�z���1�$
�zݧ��U��"	p�S�-��f���֧�Z/=����lE �H� �b-�b�D0ƸvwT���@-޵�e-s�4�C�� �����p8)'^)�G�jA�#I[��� 4X5�~C�+ޫx�؈X�C�xId��ЋM���۞��N����cm�fo�Dg$,�q�>�vu/o�S�{����^C����ts�6��J�_���~Hf|��n
L-Y����>������$UE�~ +�n�Q�0��Aw��B�g5F
0X�P�YR=�$u)��L�L����*l{Q������=�P����2`�4qv������Sݣ ���x
�������\���f�&[߄��y5� V�U��*�h���p�ڸ]e=�\�1	ˏ\Ww���}�mgv���k O�[����]�f����%�����^�w��!':��GN��3Š��_�x�`G��k��:1��`4S�P�������9��,x٦S�f�7�V0����2�]+�j���h5 à�O�RH6���j	A��_ę���s�Oȹf�$����{�������ԓ�����s`L �*�#��2:��Ѷ%�ݧU�Y���tΤ���Ѯ0�1tn#�B�.��
1�}"K*X��jmd?y�5��1�jLE&��H8�%kQ��A2�K��5���~f���[��}�(;��0q�e7>� ����_��ﾨ�,�+S:c�
��'IJ^���E.L�E`�X2�>WC.Pz󟰾,���[��������\�� PM����N�%�`�.��	B��}�@�c�x�#pg᠇�FĔ�TnД?��*�ɐ�!%",,�M(�.�⢟�$%-� 	�j��ʺ��Ϩ�=�.���(qܐ���,˹X9vK��>�Г1��õP֛*E���v �C���4�1'��b��q�)�nq.X�Ze\�tg8�gJD���_	�Z���V��hт�B��vW���x�Fʺ����B����ƕ�0W�X�؃=��C3��<w��c��U5���������'Q��l�<�2�����r2��)��8@v+�ᔹ|����"^Mf:^�P�ͺ�_��z���km�n�Q��>nDiբ��}�>(ա]�5 �^��H�6�����ܶ������c����hpl�o���8[Ϗ�ӂd��ĸ��&��8 �A���(�ײ�n�(ѻ��6^�p7�7㖵c�i�F/
�_{O���DF5�W�G=��	ju|�� .}�n0��%�)�<P8z���,	��,��X�����D�#�XH��6��	*J~�q�xoGn��/��-Z���n�A�Pb�-���d�꠯EC!�Ǽ�l-���4�'��C��S J��E����v�z:���oRB�"����9�tn����5X�%�E�
n0^[���:�<�W���#�v�]���tLSL�%��p,n6�ZώIR��h�+��R1���a��_�a>)��E��=�͹�c���Q�9s��$���W���+�<!�N�xXx�|I��`��s"m	�#���7`�*��>ǳQv���L�K��Ó#K�!��S�x�p�&�����Z�I�dŷ�̦B�'��L���w�4l$����rđ��t���-��-�4�W�e,d�6��RA�6}��%/>S�VۅN~G��T3�ᵊ��1�h�o���-�I9
+j6����w:v�4�d�M:�;��	~Ty뉺N�*���A�v���-�"�n����~�8���A�VyB��n�ؘ��^
Q�h�/�� 橬���-��n�H��pǘ��h�$�j�j�C�N�*���Qw&������<�G(�`3C����;��
��架�1�S�}��zg�F��(�<A�!�����S��?���$?L�F�op����b3��u�������vm����:4�w{�+2��#ÿ���ҝq�A��<r$9������g� v;�	�Ca�w�m��5*�D� ^g�'-�u����_��b�|S�}Ty�.X�{�jx����9��c�ŕM}�ů�w%�I&%Bmf���qIR��s�/~��8w�2�|�@�/���J+@ԐN�F)�)�0������&h���R�8����H����PU*� @�۫w���C�k������q®@���4p�5_��֠'�oT��Ɣ!9�n._�ƹ�jg&�C��:ؚ )ά(*.�H0���� }!|���B0�@�@��N�[���ⵄ�"L���5�+ޮ>�zI�΢M~p�r���aH�od�[X�O�I*jy8,��T���7(M�m�1�O�In~�\�i&��k	���W����:��eD��'�&�0��ɫ��N�E�/S�i"�x	�6r�\�Op��%�0�%L�tk�/{� ���_�׷ئ��o�;-�u�aܶ�Z3�t)ʰ��!�QP�_�b��r�������X��*���`���k�d�ڡ�*�&pNƜ6��z�&%Eg��W�XS]U��)$��|�@{I,̻]{Oǧ1�c#�-����r��zM͖��v��s1H�н�2c��'��`�q2)}�����pC�{����܏���z�a^'�0I�mb@��[�W_��+��aF�밥�>?#-E���mK�h�vF#e��o~�a>Cs��ܽ�l��q�o�m0������_�V����q��3�Q�f�#��yT�s_��o�m�5sI�-��2���q�m���5e��2\��@�(��p���[Xn�阴mbv߶�h�Τ�E)P]b�������љziz�pq�����6�Bi�T������ F�'S	w�z����I��������޼I(�T��vCcUO� S��_�u]/:"Y�{�q;��M]�q'�~Qh�~�uO���),ˀ�x}��V��x���e��J�Af��8@�<4W䅰�?>�9��յ6���� "��<Dlz�t�T�.�i%y��m!K%�����CBE��.Is�/XsSB�z�V��+�h�<�r�j:��u�b�t��UrPM盧���PUk_T�O�O~"���;��}�Q�çJ��7���XDx�H�H!� ��#ޮ�e�b�@�v��s��ݨ�2&>���Y���n�d\+��մ ¥?�-������K�a�.!��W%㉯�+ˆ&�>��:{ⅹ<l�HF{��z�U��R&��lD�C��;�[��"�ZP_�|<�>?;����4&�hr�!��m�̩I�wP,$�i|����}�)Q8k�A�}�2/#A�B&I�P���@4�ܖ�k�$�8:�2��ݕ	��k[	D#T�n���� r��j4���*�n��zu�ɮ��1N$�R���Lǘ�sP���l7v�^Z�!ۓZq��wxfeK�B8��g���&�]8�`���<j�^ ���L�JT�>3����=����:�?`I#h���}��G�'q�DU4��v|ĩ�&z���8 ��@ܖ�;����m׿
TZ5�[�Yr��]�h�B��h��3Is���O�������([Y����*�6T�-�,�-��Lt՘�����S,]�j�H#�隦I��y��:)j�j�]�t�-�D�OǄ	S �H�)��JT]�p�}SNcd8K �7�{'N0�Ebe�o3�'b<�}��6�s��'>&F&��6�b={�i?��������{lX�J�it�x�G�i�9�.���5��g�����,,�ݽ�A!�(��1�*�hos1%���˻�R�.�A�J�a��x���y�%�&�^Z�Ox5���
��|w�1� ��X=--3y�F8���m�(���:�Ŗ�A����@.RL՟�[aeਈ�tM�0Z8�̘-�2��.?VڦD/�Ԯf���.���ԭ߻
�0��SP�8{��T1���C�0E���o�jޤ�(�,-wz"�/ԛ�P�n���31$x�Q\t���$X���6�s�%�N�M{���=6KeV�/��i��۵��j�#�݇�J�����p�W � \W�]��I��o.��!-Cym�:�[[��^K������X��E��E�N?wNS�w�wz�تX�:a����O�|���A[��L����?}z��
�/OٴN]o�����j��R���ۤ=��KGV�@;�akѐ�l�`������8�So�e3l�ަ�c�ϷY��Y��o�)�$ߏ�]~`F���	S�-�P�����ig�pE�&^�ă �I��U��J�% ��g˝�+��)u݉H�KE� �;�ߎ2YB$�Q
�Z�`�Ԡ}$t6�菁e�ٰy���6�g!�*��d�NLs��� ����P�䜰A�dT����_+��|�li�GceBjy�[׏z�Ĕ��e�;gAcf��^:�>��4���I��bl
���M�cDԠ��{}�x߯�N?C��g$�u�ݟ6�^Z��a��9���w��W�fw�����1���	*6$+�o_��>�e�`�^��n����m���j)n<�@D�ʁĤ�w�^t�KOJ��~Z!�l����2�p�Q<wB�K�cNG詎���\`��������u���W7=�8�03��~�a���4�R-�Qv;�,�B�%�WAIʔ�k�a|:k(���s�И�Ҁ.�m��[u�1�����.>|�o�;x�z�}�r�t B�D�R���.�t6m2ߘ/̶r�t�X�<�O��:�*�V��Ư9�1���|8�i �����%_�#z?1�D����!�m�y�d���&����w�T-�wHN1�Yk��>�~��e��í����R͗�K��0�ж��I���O)�/+!��T}-��,�l�4����"ɸ���bG^G�X[���E%�VR�� w�9�T�֧�z�D�;�Jq�;CejGh��G�8��L?�f�:�PJ�{T�C�9r�C5�9qy1uyϔf�x�T�9$���27�����W��K}BDTq"�Wt���%"�4.]jb5g�˘��s��J?ݱ�(���V8�_J��w���!�	�����D�	�`�c�'KkԞ��?gJq��{�8��\ �P�&*�m������g�B�^m/AyW�ӈ�2K)3E��m�	Zb�ao�a�P�^�np@�����I��M늾�I��s̊Z���=�"���8�D��O"x�?���]tk_�`Z٘^�@���"F�&Q*����슅)q� �6�^)�x���s<�Z��Ek��0�o����9���	�������񆏴bq���w;�I1�I�Rm�&�7����j�X�u�J��F�����ݝ:l-�l����a�@��(ޠ�>�n��B��*�{�v�8�s�<�qz!n�Ҷ=�q���f�T�m�ܽO�_;��"7g���.E��Vհ�Dq4��\���Pt�b���L� ǟ����$�	L/�+&O�:7�5�ر�N���\r	��x�:4B�7�l$+g{Ex,l��2O��'7����2�8���dv㸽}-^Yŗ��y�\��%�f�����7����AD�h��+����R�����s��FI��̐X^���4e&�����2�u7�ԛ�'
c�ATj��e:�$.����R��;3Zzr}� �M��I__X�2�ǝ�9����K�Dd��A�sP�Q��D�V����t=+3�R���7MEn���O����z����{��K&�;iI��r��@��7ʹ�~�u?�D0-��_�4�l$:6� ���a�`ba�해rB���������l5���W�}ٴ�%����K >tF��W�JgvE����,&�a%��Y0�����L
vԇJ�龒`c�$�2���x=�Vv�L��x��i��?̲O�^b}�Ѷ�D�i�����	E?��$�����uj�2��	Fyj��2�'��=l�,�}g�� "��s������p�<��}pa%�\G����ᚷ�+��Fj�E[U�=ih��;7&�?�3�y���!��3`Z���� 1
���Zvw��q[��S�{з��6������� ~Ր%���Yn�Ct;�|�U�~�6�_e� @�� j�ɒa�VVBb�;b�Ј}=n�BN��aL2�j��-�ۙmEV>�A��`	�UN �ʌ�m��$��T��ȿ��&�^<O����]�~�	���*Cʮ_��[$�����\�`ȹ����֏�l轴&�;k&%��8b���)��c5�өk?���x2 �' �w�c6C��8��Ȳ�\ޖ�DˬN�E9� Σ�Y-aczgز?���MS"�V�5�[��}W"d��Dy'� 
x=�u��~}�R����>[.���6�j���W��\@�!�HEa�yB�]DQ`k�#hⓡ��;�k?Q�v���p�`#;��@����|��N�GaI��-ù|��P����`*�3\+��H�ڂP�B�W�*������x�]�婈�6K�60���X�W����D���3m�e8���C$�k���o���W�P�jn�.�-l��2QdpI��.h�gv���TZ��ͬ
4�O���k� ��Q�De�Vm�EW�����d��L<��K��>N�A����RU定&�4��bğ���۠��v��-�\��#���i�9q�y�7�,��*��߆���� t��t���2��c���sI8�?�m�48+G�<���o go�d�|���>���WR�F�CrDr4�2B5�0A��h1esЯ�?7_q^�������VĬY�L��@v�jq�-�Y�_��jz)ТU�&�*�5����ߔj�D�ж����I
�)��]ZSԩhb����tm Be�X�w����h2���A�?��}�Y�3y_�֏������x��<o%&K)�f�P2&����欆���އ��=[W�R谘ށ�o{^���E?��B.�4f�2��z���ɓ�.+!cU���K��X�/��3D��F�S��U��n��U�ͱ)l���9Ywf��TNfg��{Z�+�ug��[Yt��I)����r+��SNT�zcǞ�ݸ�B�8Xn��v#rhŠ�i<m��B���-���Ź�F_��<=0�ݵ�ɦ�b̻�.#�c������+�6U?!�P�H��(�S������O;ʏ�.T��v.�xL�_���eb1�g��ɛ+�%�	 ���	���e�<?K�I��R�-���������n2��>��'�tk�sPWᜫP�Q�=��<z�;��!.�N�U��<�Kw��j��/��G�iޣ��G�H�K��t�����|l;3Ӆ�O������窭�Y1����Yt�
a"���Q�am���Yk/��oC������A��3IBa�ݷ=��t��J,�+���ے�|�n����)HSQ#��j�^ro�ձ�AF�|<(�Q2گW���(,&nJ�Т>	�q�l�� �; �Yfp�!���<%�������c��ie/6|�-�ieOe�cv��"�Swk��>C�	P�0�`V|ru���mU�C�֛WUvkg�x���h���[q��1"�
�ӟ&W�tW�&����;��/�ȴ�R*��>�W�C�m/��F��e��/�;Q�T3��1��~SU�R��t���F�D����Mwq86w��7�����cI�t��+���(9����wW
r�x���<�X��3�l�-��d����|#���"w.ς��Z%������|�7�'�����Wz���f�����?7;�&�y9сvx�7@'�{��H��n�P�y��~��d$�j�#~
F�ыZ[��:�7�+W��������j�H�ZOq4tZ����)G7�@+;Vt�M���`;h[���M�6D�1�e&����(��2�l�'$�z��,��b����;�Y��Ԍh�O�~W���̤a�ލ����d�I�M�X���䵂�0V��xΥߣMaM�0%�lT�N%�k4��fh���0��d6ET����2�\��N���ȶ�D	�^�v�WlI��ݢ-������?��Bi��F�OK�Iga�Ro�*�D_h
<5قK�Z��D{�ܚ��J�Q����8AK��)�����/������o�a�S�1�D�R�L�aSZ����ex�0�u�H'�l�=��n:��d���1�CF$����VSѵqc�2b�$=��m��z2,�;?��2E�S>�c�D�_�Bj��s4���������݇�]ӏ�)�x2�y*�J�Yy0���=�%Hb)�b�����h��y�X�ͱ�r��:|b� ��Gq�H)J.��U�y��*~�[B>W���h�X6�+��|�)k��E= s:�pӑ���c�W��9���%�Q:���ܧ�˃���G� ���H���H˖��\$�˞%!@��G@ЉJ�)H%�I僱�W�Ba�� �̈������}rC�Wڞ��'��ǡ���#/��{��፾��@�a�B��o��P��d�v��z�V��z��-"b����/�T���:�\�6<iƘ���q�0;�²S��'�-:��E���Tu�,���R�G��**���Kv�%<�ֻ4�*J�te���^������$`^��2|C�� _��&h� Y�������c\W��;��_�\((9�\�}r�욕%���2w���3��m*J�h�� +�I�|�~d�]tX�n������B�%���nM��:��"P�<�E�����=�V�/WK3�O8T�����V��J�dt�?����d?+�i�b	#��KU�Hzl!�J��R2�������U �6�"��� �/�Y�fw���9g�lGFX{�@v*"	P�l"��c�G���W-֕�4EN;�$w���@P�kv6	�GkvD#>$�zdn0��^|�}D��.�ά�����(\�r	�[�-�W޲���#ń�����3�ඉ��x[���]�^h�+9L��P��;�w��?�Z<ܟ}�I�qL�e|:DO���8 ��GH��D���Ќʇ8[Q����r_��c�RX��&C�����l#՗�_3ez��n5���ɽ�g!M?�i���*ty(���3�]1�D3_<2��o��cRH
e�����;�QSCࣞXKl<�1�؃�V��xaS�r�>��c�/��h&��&��ߵMѻ����r�ppk�����.���)�0)
h�� g�k�F����pq�F*�F��kFw�80�[)�'�0,{�`B�Cb�I�Z޾�z�8r�@ׅflg����]Q%��h�a�`n�aTx�|�;)�S;5�QH@���C�Ȟ���_�=��cl�(2$�����ea~����<�0����1u�^�_����Av\ C9UT��d��:��x�ϵ�p���}��r� Î�>�
0L�����K��b#�����ǳ����\u�b$&w[)V���Sa�Vf`f����\���#��OG,�o|�uL��:��B��Ϋ�Z>��U�
��Ik��ѮiQ����Fp��>���f�rQ��=R�j���b��
C�5�R��i����HE�<���BG(�(��4y���0�U�/i'�A�zl
�RЬ�-��:t���"��0�pK��@ڴ�M��V.";|W�1��ea���;Q7�:����I9r�ւ^:c�s4�	�k�o�WONhho��! CοV6�!�Owj|>����H	Aʤ^&���2 &��Tp߆���uy1u7bGs%S�k���g�:c��ɵw1v���:���`��Z�I�)�p����ט�F���^�I�]w��?�Qc�4P�Y˓���/ve?`�� ̉2 ���8a�s)`�MS�D�x��g��������c�W����m�[W�p�aƁ ұ/h{@�@|g���h��kb��{.��^��;����+��c�Y�&��$Q���G�e�u8�K�oJ�~���`��H�Z��e��;��-16�m�y����F�W��`P�x�Zb�w�'&ɚ�j]��-GP ����f��i��Ŗ��k\�pQ��:8+˝�h4'G�*�t٦0��K�H���g�Jr�y&S/����<#�+��+EC���V +��.�
xZH�6��e����ݍё��rQ��E��_9<�>�	@�d_�bE��qW���%}�W�HtV&����)Imz��ܥ$x�x��I�G����熕Y�L9<-���W4|:)r��$��}f��ę�Kك����ȷ��	���Heɨp��}�M6��0|OkH�4��&����|nw_l��'�(&�o�~S@ٯ̙"����YV�v�h�D\쐶�i���W]fޭɽ#,�%��$�/.j1�5/� �)����$h��W��r��f@�WV����6B�to���+o�ǯoix�����%|,��ktc�Ѝs�'���wqJ;�\��6�us@����ͩ,wb��@��&�d3�Q�����Q���bc��<��ࢢ����[?H�	5=�T@|�Qg���<@�~�^��%���I�p�/im��\���";}yՊ	�;W�����9㞉��*_��"*ݳ�׋��yQ�"/P���������\���`(��[�R��?���2b�Z^�6��铅��퀱�bb�B��QކxV]�B�N���;�I��8�U�d��q�(xwۃA������7.sR>G�A�~ğ>Z�niM!ڜC.Bqpՠ�ߏ �^[�+U
�S �@<��$�L{������2�2$�y��4�&�A���F���r
�j��WO4�=�+�!]��r��↍�]tѼ�E]!Ey��t(4<���UO�?�K�� ���Q�>�	�6�*[�;T���l�ᳮ�U�1�1���D�V���ń��O̗QU�t�j�?����D�#�Ѧ����p;/"b�U�Khd{�f��ٞP����(C4/���<�:��~K'9�?,���������o��cB#reR����Q�B����
I]����2��"n�4�I^=>�PC����y65������Ǟ4��o��$���c�T��Џ:���fq?$h�(�'D�I��0��3�^�+�]��������E���񥉧��,� ~6�ڴॸ ����%�Bm�\���*<������W徝�x�ʏJ7!q�K.[��^�d�4.���/��!��
�>Y�lά�Ʃ�1"����m�%w$��lxɔ�Z���f+ic�����	��29�����%���<YD~���!t�=�$�)�Z9��H�z��� G:�y�Ɨ��6�9lh/c���-uΧ�G��i*�'��sU�]���,�%�[��Ձ,��0�2�5���{SX7EGG�����`�㖛Oha�}E�����j�%�4 C����}2�7�n-�7�=��X��<@����%�6V��c����A�����ט���& ]O3�p�Bx�MG�w���k%�f�i���Q�q	<�1!2���d�׌C-�`��ʞ�4� �h��}��oA�++zAAҟ"�f��Y
�����+<��Ή�ŀ����w��^���x� X/���v�X2"�sԌ�G���A�r���)G6EJ0��K��������Q#� ;`=:���]u��p�X���`�M��Q��^B���(�?��ﳬ�CI��ys`JyÉ5D�tfInW1�nw�~�R�;wD$�k�5�v�P�$�_����c�cp�����%|C�r�[0l�X*ĮF	q���5�v{F�b4F��`,s䴏��f�.N��Ie��:���|������D�M��(��3�+,���8�f�P��~A���3��Ї��wqZotN��f6�I�-�`�B����Z�]�m`�0�&2���^������c�.�3\v�7T�ؐ�FU�R�nARmT}��zD���L	|"JT�e�Pϙ�ϲ��?o����fB��ˑ��WFt�4�:���"��N�7��tF���M�+f�*�� �ɜ��P$�f��M�ѕ���	X�Xt�/���E&xxS��P���uz��m�X�O�:S��׊n�v��\� 5)ğ�z���%z��-/M\+ܚF�'�	x[��r�z��$��K�
��g�E�!c��%?t����� ���SdsE
�2��DW/��������e��dz��*$�?�3!�d�����.���zKmIX�ļ��3ѩ8���î�'�L٠�P�8���g<	�ɥ�bS���Z����E3�+a�6�ei�^��*]�ا�A	�E��=�����	1CHѩ�~(�|^Fk�y%.��Q�`|5���*G�v�(��e�2��(���h�2}X�^�?��<� sR�-`sy/r��W�2��G���i��\K��f���6�1Fm������p�N�Y.-��[�I&84�a�}3���@��Gl��uVmв�2�
�Y�5hb���T���Qu�!��e`"�{��{�8���)��'�;�s���M�!z����;�]���N�@Q�|��׺U��l^6�Z0>�h�P��� g�D+N�a�hV΃��(^�E�HS>�&�]��.���9�h�Cԇ�3�#Ե�G�I䠡�@�W��M���=��mi;��s��u��3# ���Ҫ���;a8G�h>����毉y�h�'A1��eV�r��
����*�o���
�4��}�V�r����UK$�/ܚ�w>	�jo����?��3u�N4>�]'��`�PyA�T�"�]Ƽ>�m��"�CN9W�4��%[=�7�k�U2HylPP>�:�惑vή���V�:��57����/x�w�V���Q��M�vVm��uGN��D��痲f�bl Mo��(�̱�㍲̓C��@�kv�3��~gX��f�pH[�f\m�>���gQ)�S+���;��,������<n�v�x�-��	h��&u���J�҃>�c��b3F��}�κ\p�4F.���O���IX
�P�Mj�ط+K�V��������x4�lX6�Qu	/ޗC*�zMm^O|Bݭ�iB��`��t5j^w�u���l�jܔv��|]���nnl���Aa��{��$Ѕd�<.Crm�'-�m�d���ֵ��AU���eX�w�Z.�X�T�u�Y`�UgZ�Z�1��6/�B�"�� ��>SΈ�:���
�p�ǩ���-����^����/ܯ�Y暳�@bt`��S��
�%�;-s��-�2��`��ղ�ns��r\�D��}����t�Ǻ->��;���<���p�Y�ǣ���=�z��7I4�AMb9�EB�[��B��$s��1�۩�U�$a������x��,$�O�{��Pu���Z9�f��9�$���ˌ���!��XBD��O��% �+v���7�z �Թ-�I���ز� ����|l{���A[�q����.@ǡ4�9��xg2'�Ȑ�PI\�x䕉�.�J�@��[�r:�<���h6
����sJ�J��+ռ��m��3?db�M��y(�{y����tͥGIzz{"H�i?:��Zo|<�y�eṰlY8]�>�شPJ����z3�6!U�1��0����\�=ϥH��+:2S�N �]&V����>�| zל	ӞK[�+��1�-�& 7�hL����3\�ޛ[�]=ϕ8�x��ϋ�k��UL�t�#f��)F�����N!J�ѓ�s�,SPd���W��%��x��^���K=5H���i����˰�Y!����l�d�R�҃JRkő�?u��-�*��aş�A�ǁ�ɑ}�x� �4��+χ.BP�� �,M�rDf��_�s���K
���R�f@�y����3�p���n&h���_�S�5�m��E�#S�Ҽ ����<)Z�1�@դ|���{+��<H���M�7x�|o���a����uHΛ�I�>��L�L]���������Y	�j�@�n���x�Zp`�a�T붓����c��}�����������@6���\ޖ�~=S��V Ť��=/(�~T�n�(qSڷ�U��A��&"����d���u[��o�󐮉'2�|�YO�Q	�O#$S�n?�z�{'f������W�2�gW=�ߙ��5����84�;_�Ϻ��p�?�Xv/\_2�t�%Ŏ������ԥF�	η ��V�P �_U���pJR	�l�>�i-�(�D|��H�Y?��5�CI���`���H���X��1�H�=Q.xی^v*�Ғ~�G��AZ���L�u��5��!��K"L�خg>���/�8�ͅ�SuEiж0�ȅ���.oD-Z+�|�3_���w�ۥ�ď<I9{�k��(GŎa��wp�6�ܓ�If*�$�	�d�7*��j��T�$�BȄx�جt;L
����nne,**Y���v�y��LV`��W��ѻ�^�W�ɹ}��`i�c W��j3:��� FM�e�`�@e��P՗*�u�4qH,�q�-L��o�x��H�B��k��P�s����?D�O<	�9K�������J��~�)8��rE�;���Z]�7P�����W�o�u�u�����Ȃ�i�8IkǶG�0�c� l���+))���������ƨS�Z3�n��J"`��wa27Hi�2��*۱���i2�nsC��0�{I
�̝����_M�����i,��)i����f�_:XX����ɉ]����~���ݯ�l9RT,�3�)B��~\�¹Y}!
�֜AQ����6^BPL�
����5�r� ���cxZ�D��A�TI��m2a�-BBg��4̖�(����/>**�%R�^�B�s�p� h���y�p�Ss�Ρ^�b39�#W��5aQ�y!�}U܃�.��WjB�=u�ߴ���x��F[W��>d�o'@����&�����F��ٽ�`q�`փ�vU��|�X3�	��_ ���8���eoK���C{h��$I��o륎�_�޸%��V��*�fAd(Xł!E�l��%.{�5+/Bj5��0�8B��9�H 	�1���4ǉ�2��f�"��ނ���/�@9�u��D�"� d�m�Hռc9�/mЄ�Bů�$�v%\�7�. �l7��X���?��3̝�Z=u�I=I�3#����Ha�(��v�#BA���\�]�^��gEp����]"�t�b�e��^�J���B��"��
"�}#< ����+����9��_DJS��h(�����.l~��r�fr F�E��"z%��~�v�F$��vr�:@�����,�(�6�D�zfl�dTU����~���^w*i�M��e����5rׁ��\œ��ZG�=��JN6�5�(���P��&����4d���"��qN� �K����?��e<Gl7�k �_i]��G]��=����[��cΦ�&�#�"����E��0��{U�L �Aۚ�R��*?v/�9FT_W������3u�^�҈�p?�.���^��J�nI��:q!1[G��ƯX���]��Nh��du�m�oM�L_m����Xxc� ܈	c|�i\�6f�=������Z,q����<2�\�KR���_P3���R&vMW��E�Ѽ�<��?��r�[�Y��^ę��y�޿ET�Xjħ:�7�E
r����*�z���Iu}6�����'����$=���Uǆz��L�M1�i���ϫi��!ME�ٿ
ʍ�ZN�����W�o$�ݦ�Y�`|3�^�C�,=K����^,6�B�!��4��j��b*g�����q �e����o��o��x$�R4M)�e��]� ɰAl�T9p�p���/�ͩҍ4a�~�2˿�"&�`��r��0Ǔ58���ɥfN0���M&�������1��԰����'V����n����[�NI�M��ѰE&qb��})�3l'e�Dc�7*�r�Jf"m\�lq�a�T1��f=a�	^3��uzLǖG��|�@ǎi4"~:���]mQO3=_�չ�3����TM����JBA0��Ǹ�&�[h�&%\�|D��̖)���F�|)u�0pl��(�#?tÝ0|G�V��C��Y,ǰ?e<�!�����6R��R�̩ y}�<Ҫ�.�A�d��	��B����pD�{����M+�����mq����i���6c�X������Nʼ���'�	�Q�}	ƙ|z�����ژR�N@�57V�,
ΣS�ې�3鹴���MJ�������t���U�%BV�ˑ����wkvy�3v�1�]�G�A��y���YʥE�7N�YkZS��ǿq�"5�L������9��|W��*.�����7-l���}�yNy{u�(`�G�=�f?��0B�>+�tL�B��`3��A��' j{*���~�'&�ۜT�:����)�Jb�F�+�`�<g-���cD+�����v�4����/ whOxǉ#a]㰍���-zH�#��VƉ��.�
W ��a��h�XT��\�1~Do�}�1���|�'�����A�@���$�Q��	_ߒ�^)8ȁN��ὑq{so��|mȅoY�m�\�w�CM���(�D�~����6�t�E�{�׫�#��?C��
z����j'z~��5{��	FgC�?^8V��;_��Ob֛"2Rg�WDʴ y�p�9���u��52!�&��9=1�|�;�vL̐y�$)�bz�Х��_�(p
8r	��-���M?�g�ss�|�f(�-�Wf(�@A|]M
Kr�̊/R;Ԯ�'���숚%���ǺX����M:�����`I��>��	��G�ߗ-�1C8Ħ��������]W�;��O^�bWS�D�o7����R��� sH�:T$é��af�tL�Չ���TȉDҞ�iI�>���l�k!N1��d��j:Ё�l�qڈ����쓃��� ��J�=��6츒�RV��Tm���.����0�H�Z� k!=���H$���c��X[��Y9k��}����υf�ҳ�����bd�%�M`�$��2��{P�H�-����SҀ �0�a���������r���h�O�g�W�z�	�W�]%�-��.d�w*ΐ~EI�ʤ�O�kem� C�K���U��h���/�g��a�X�2�:O�K|wz:3�G�g��y�ru�MW��E�R�]XV�-��b铧$Oׄ���2��y�(��%	�Ӧ6�$����#��=�0���'y��S��`Q���t\8���[���77D�3pk�j��'�V�����E
����]LzQ���-�^9ox|��dm�8k����y\�.G��r���y�A4߹/��
䧵KZ ���ʯB��9C4B�h��E���b�����`I��z����:ZVp��/RԜ�܀˿�5��[D��C�������|J�-��ߍ�Q�˭��y�.z�*>��>��9]-V��9H%l��V�̴�}|<��Q/�w"�A�o�'>ƛF�hHe1="8��X�VT��z&�@P��?wR�$kח�ȷ����F�T����^to�5:�Z=~h�I�c̹̅�wfM��UlC���6�j ��J�_Zד7�'��{P��O~E��~�Hq�v�P;J��9�*�xshI�k���U��ݦ��>�nH�a1�E��@+p�m�aԡ{�1 �ats�@�e����<�k��&���|�O$�?D
"rGy��r�7D|4љ%Ê{����wZ	������I�M���G$<������e� >4^����t1�4��y(�{)�n������7%�=�HV��8�����A��=�J�:֟L�'��ߥJ"�Zս�2_0��!�^z��Q�c?"�9[�rQ�jƝE�航����G��:6�t��a����
�7K8�k ��+h	_9Z �,��oS?+~�"Y��H��iM<�W���L�#d���Kͧ�8{��4���4�#g����tŰQ2�l���S���џ��B���1���?�ީQ��;�i�TG�w,�-8B���d6��B��� ���:G�&2��l��X�E��ybq�3�w��^D3����>U�C�QA��UƢ
�/a�%q�5P�kI�h�_���d0�MD�#Ol�kjVF~Ѝ�-M\�7[�<����G��퀂e��[�2�$V8�T��W�C���f𲍦]�\�.��j���x�N#7[��%K��H�����i�����ߌ{gL%�_x�Zz��;�;��?^�p^0E���6��T��2��:��{�wz��av�����Q���Πl�m�����u��J������e�N@odO`��+�͓�+:�&���2g��%�J޾,m�Mw\q��]���{y2_@�SY#��$���#�m�1J��Y�֖/p�<hE�E/q\���d6��/Ã= �
v0L�C��`:��%�����#rL(7w��mԵ������R��N��8,M��ݘ�LK��)��ѱ�P�pF�*�V#[n��	@��D���9Q����(�l��}AZ��˷׃�����iˏ^�v�6 3���rp��r#_V�
PleM�$�{ct��'`u��T<f��T2���l�\\*%��q�bq��F�YE�'��5���K�=g_�>�Z��;-^���ߛ�VE��$��DqÂhc�k�^t]+�7�iL`�������֯����\1-�f����Q��aq'JZ�����G�n�]&�_lb%!P���ͪqܢ�,�O�����6��
=�8E���.8MUP~Y^�w�'��xF53�ZH����%��y:��C����^��������͟
�2v�� �	'�M�/g�N�����.rᰭs�e��ĩ�Ff�p�\��Nt���1On [���G�79Fn0/�g*���^�	�.
��{dM♹�	b.��8 cYQa{�P47��,,WŠcs�ޟr6!���H��f[�r���>$1K+�>�:A̶�睗Xy-J�@8�Q�>�.Oǻ����r���dN�
�B�B q�E�5m�N������K�ßXb�pl|k��?a�):b��h��|:z��Kb�ف����qPZ$��=]?�hm�F�<ͩt���Mp�nn�� ,?�r��:��@S�V�������KŹGUF7TTΥ$x�:ܘ9�k��t�����6�7�d`�'K��:l~�����>I3�Q��X�I6Qq�^ӿ�8�`(9
@����%�A�! �����f�;R�F��[R�>��b8Ah>��=m�X9�d.����+�+og㏛����J-	�пM^B����aIl�R'Y�+O� :�5n)H���*���닖w�s�TS�r�rf������궄2� ݭ(�!k�~��>+��� `߷�������'Z	��a�R'uq�C�F$v�+���I<�n������`�m�F�K{-������7����9��K- �������b;��*�6���-�n�y84-8�*k���֘;�ހ˾p~�clfm���Av�)�m4�;����ٺ5�#����dاGi��wF��OD6���q�B��c��ox8���[=��b+�Ȫ�􄈏�v	s�@<9<|��KH��7P��K��k�e	�<�z�#kK��ۈ�\���|�8�g[�!>9�TO�����~��\�2��������>S�A���d �!3ط:�Bv�}pwEԐ�l��s��Rn�ga��9�9]%re/��>do��d@^��2 �1�G�y(�]�"nM"vCP���-��j����I��� ��B��E��z+���s*l�_���7)�X���tHU�^7�x�8�Ge�������Y��#նU�/:?��� v�,���`볍OaQ4k���U[���&�N���r�j4o�=A�7&�M���1&0tbnC��P���3�W��L�dI��ة	�+0=-��?|!��d��9	�:��o+����|�2yЌ8�1VSnB���	���j;�!��`�荭��+s#v���,��(�S��#D%��0g�9�\���ق�+�уa١#�;�����Οa�D�˺���w�˭�t��=�'l���2\;���Ҋ���pk�A�<��IOб���`��xֈ��.��IPq��U�>%����o��ﶥ!�� v�~X�\Z�
8bg�Q��L��~+��$k�h� b
 4��X�fU���79��l�GS!�D�%��,��Uas�"P,
q4H����l���N�s���z.�s�P�GQ[5Ti9�؃�2͢@��=�hT"Xvb���pv���{$�<��"K���jXV�m��NS�p�=@�F�I����0���s�d�eB��AE�_su�������V���O͡	�jJ�U��=�fCf��.�F��Y�l?E��)���r�*��Xt�&ZT�I�����G�~Q���*��S�7Zre��L���w٤6fgͿeO��js)���} i,xj9�-ϭ��_+!<!-p^�~��$a�9�UGy7�Ci䵿�H$�;E�K�j��+U�r�ƛma�Dk�1��4(���B����ډ\������i�ı3�'��O��֓\��=-��fO�� ��x��e�^S�o�~PE��v|L�4�Ϊ���))z���<+'z)��¤tivQ�r��G�C=a��g4Ga���x��IM�U�n5�D��_4r%v-�|R�{�[�^����;�L�����e�����~�a(!/�Z��?^qU��-?�\ə�/��t�W�Ubq�<��셕2�%����ѵ�2L�Q���T�o�)IYV����=X�h���d�7��5Ċ��S��w�MM���I�o��r;/~8 bU��n��>o�����8��-��S�R};b�7�@!�Hk��9s�׳�^*q�Jr�W*�H�
�:��q���F��2���ؐ[���1/`��K�|��V�9vOݗ\�S����'$u����
�&���߼(��6<5D̪�t2п�s��Py0A����E3� <j��Ф�8>����`����E,py�ؼ^1�f�-��(�\#��)����[��V ���ىi����u"~ۉ��Nǭ��A�� k�k&Q����o-�@��e�T[B`�COV�']��p��������^�m�8��1���g�5�:-����%�U�	3	��vi؍ ��k��4���Å�V=�R�y�a�"���`�jQ�&��"���v����gh��勅Ld��^�t�)&��ؕd2�p�||WJ�0Op�p�C�X�i��҇&/A�ިZ �#��1q���혴sk�uݺ�Ƌ��B#k��y�!X�Π�����x��k&��&�v�I���� �A蜰���;�u7d�,��������o˘\tߍW=�"��>̲�u������,�^��LXN��G��"�k�O���Ϳ��UI�0JErZoՠ�3%4t�"��9s�F�c�O&C��KH(?5f K�:����R[��EqK(��5��iNU[���H�=.No��3Bf�+*z���2g���F����X����R��ȢA���Ϣ-�D�׶��3�0����
����>�"��I�N5�Q���!�{χ'F�MN?l9D�45C������dEƅ~��|�6�Oq��43�ȻW��gų�l\�H	;�s>�'�t�F� kN�}K�E�K��ޔ����}`�si`�H>��JP|R�~ ��@��9[4�������bQ�V0'����*��<,~�^{j��Ec�8R��y"���}�?a�t⼽�W(��M����@�nz)͎z��n͟U�qxȼ"��Ti��t���j�DOT!��P�렍*�xY����{���$���.�����S,SB�8Ԡ\�]x�j���v��U�7�/W*]'�@�i�3��
���,�<^	8��;�ov����	�kX��l_�������a>� gԄ{:Z�J���iѡ��qd�p�H��uV)���v�H,-����߉`��;*����^��ע��,_�.�d�ȸ�88c�ne!������4m��/��� C��;��͕.�8��kD����p+8�$���T��\]����*�: j�d�b�n,�)m5~Ur�T��D�O���F�;�}ḛ�������D����$�ho�B�+���#��?�$��1@|�G\�f��T��) 43��9UEO�01�#�d(ȏ9�"���(Ti��}�|��r���<��Jjܨ|�����dB�PZ���P��K� G�V�9nBA7�DP�̍���2��{З���Qa_�<�z7ˎ�R|�9�&�m}��p�
�A�du#��D�\��׌M�5�.tr�6	I��b��渠F��D�"�����݃~t��%���8U��}��z�$z�j�>m�ü���|��6�Gh`�&Mg$UB'�����@:�,ź�W^��G�L�~�Lc��W\����c.6�K4��v`lz��{Xb �=-R,&�-����ңV�V�[�ä�v���;�X�-��!4 (-<�ް@�s�̏ 6'���"�(#���~��;!���s��A���}��ȟ�<����Vд�Ζmٯ2��V/(q����f �b�nv�?�I��o�FZ�=<�Y~�<�V<o�� ��Mz<�'ԫ����� Wq"-�M����T{��<ę	�?
e��T�"���%�i|-G+6��/�C��#aO�5*ücF,��S� e~��4׫����p�k��l�N|�b� SSc�V��;x�}�02������>��V
�^
�$oI<�x���$�� ��h��4��V7uF���&/qr�Ӛ�
W����|��$z�*�oș����`��h���v�(1�t��o����6��|&�Ym��Q�~���P��='(j�~ڊ�����p�ǎ��+�^�X�Pq��^,���]�Ry:�͙a�h�zӦ�Y�o�+Ƶn�D��/��J�������2�k	'^?���U��V�O)ӏVV�S0Wl�R�m0�7-�5mC%��sz���[R���5�P6�c9�����o�]�M��J Cs��ٍZ���s�k�'��>n��JD�j�[�	`@��5�� (�[@�ܹt@ju4Қ�+�BHY�`�}�/�J��m�N�I��ɠ�3��so�s��+�ȥ��?�Dn�C#�6��􀢘Ȧj!��9t����!��0�	��V�|҃H�h�Ꜹ�����!���|N��A�8?�\�=�S��[�1�W�Xsl`p���Svr�D�\�,��m8�2�N�}��H~q�E>�Gд��|���Bn�W@�52��/ފ�n5z�ph�Հ�(��l�4��U���*����Q�`�]�fƷlT�է�U�t��/L���bTi?�O�t�1]��٤�A�s?�CO�BE4�젆y�(���B|��vĻ&	U.���a��D��:��U�^+�Vq4�$��+��nw�ڈKj�#Z�#�&0�}.�K�o�
>8/o�Y�"�bG+�H��S�3��o��n_
��ž{�Y �x��{նt���j�QOw������7�uO=Í2ޡ�}�1M����WhԻˑ`�5$�}�Jv�����H#�_׬+c@��O�ёKuӜLa@t+Ӽy��5��7I�5��Λ����h��Bth��w*H�I�|�)�Qj�$4�K�&�Ԛ�G.9�S��.H�tB�E�����-3:�Z�s���`)�";�=��u��S\�c���x�A3��	@���\-����CPB/����	t��Z� �d@8�O�]뻭l�B��({��^��$R̕Fʇ���:���t�I����R�]HD��g?oa3���L,Ȧ��_�e�9&����h�X�8.�)��~<Aӑ�e�)+��O�q��ꐹ�y�D���O���b؅��ZH?`'���B��t4� ���u�U�f/X����_-�S	�=�6�
@��rU�}�����ɭ��Y%[��^�������,�̯#�E������.c�OI7�K�|�xl���� ��y�K�����Q�u);:�g�b���o%ML;���^��=��^��ؑۮ��]�����4m�c``Nj��9�i0�C���\eܑ�5���F/+vdF��(����ݖ��4���8��+�='��*�c2y�Ŧ<�&��B��>g
0B��,�sw�D��L��I	��M� [ 7:��ka��m��{9i Z!&���_����@,�	��m�5菭����� ��E�m�3nj/�$`�)�NYF;��y 6�8�\ �(���f}��3�Qv<��q� ��>^���y�`�ʡڠ5��ā���:�no�阝J�ɇ����X�$.���^t�]Ǥf{eHtM�h�����B�rݼ`���M_�}���~�5���G�����i p)5�f10�a�b����<���������S��V�o���@a���\77�������2{[�7z^�Ao�7�3��X&3� �Q>\�7�iT%�U�ݡ�Q5D{�gHR���1R�;T��nl�^6�%L����w	yaz�ÿd<��N�"�To�Rt����X������~*��#˵i��m!aƊȦ�t�YL�	g���
��B��k[p@�_%�Ȝe��@*�q�����N���ƈ�&D�,#Հ9
s��=���$dD��"'�ҧ-�'<eU��_�V�s̓���-���B�N�����Q����(�9:��ϿO��I�*���1�M�˂@�8�m�n`�|%�.Պ�=s�@j�O�W(��UU�c"YQ+,8���	M��ц�˿�3A���Ɏ�>�mo�4 �xF�����0R�I�����t���V��b��8�a[
'�,�d�F�o\����8y�����[��Q(٨9�����6@�]��x���G�A����Ɍh����g�m�5�R+�&w�r���v�"�W�0��J>H��Xc��,�O�3;��Ѱ_i��hJ�(,�����=�DV��j�f|�~Ɓ�;�
PpBe�X�4�d��m�D��3;�!#��V�#Ӈ�EM69��ɡM9�F�s�������{�a�������Z��eO](d��}1��Fg!��������8�+"q���'��MՔ�(Zz���Y�.�l-��fQ�hI�<n�!�َJ����K�m1��g�{]B������u xQ��ޘ���@o$�-NC�����6<J��>����)sc��vYjC�`���ɿ~,0����\��'	-�h��wW�Չ��_�uF��A���I{�fT����&�J ;�:-�N��<�����{,HF�u�����T^�Ή�1�j�U%�][5��KhI�Q�K��<��[�sђ�]���!!�Xa��1~69�j�O��E�feC2=�R�,�S �wE-�`9zq���*��h3���w����\�m ��{�O��ΐ���*��	X��>�̓P����D�����	��a+���њ��[=O����x�Ҡ�P:�:e�z c\��4�X�[\��h0���h�El�}G������K�ݶjLD��������R�x?��[	b�0�޻�����a�2�A�A�I��6�Ts�6CM�;o�o��|*h��~�=��*7�>��o0tT���96�{��bkaMʋ;��>��7��iP���c��y�CѠr�?P]�<׈�R�,s���&���+Ȝ���CK��,�����Yگ�y�	��`�"DV�k���V�Ѓp�#@*m�$H�JA��B|�[ �@,cW0	�q=�"��r���BN�#�fL�b�G؅���x�+[s�R��9B,�sӲ���I�"�t{D�L��3�J/�.��GƗ�����!��$�E���v�bI�(9����b�YT��s3��5��.q�� @�C�]�Q��z�.8&�?9f�,��|w&[��
D+��'�!��˯��Y[�}b���ߞM䲕xb]O���]y�s��[:n�Ԕ��f��4jH(�^IK�x��&��oDE[��{I��m�	9�f��ܫ���S�>�o5��j�8";����E�`>^�ʲ��-�&b��sbf�����������}4r��OYP�%�]cC&1�Xuf�}�I0�����E�[�0�BN���(уxӌ���sɴ���9&��oH]⿡��������<�m��dc�%�Bl� 'T`::���m	�-u�3�sNZ�5𔕒��r��h�Z�Ե;��񿨀Q.U�\ ��h�T}x��v�lDM'wRu���v��Xb?(LHrN�C���U�}��Y���/�'�Iiz	��;Pм|��Ӛ�������p[#W��R�L����̇�Un��Β�_�mqD-��/X9uzeRGT�G�n��|�Fx�[�N�=��r_˘��}:w=�%�,�W0K�G�N�O�"9 )߽4�J}x{�r{ Nc̐�SW�G�y��yzo�a���630Y�Ď?�`�,C�^C�Ș|jЗ��(�e�~�a�=Y�kh`0q�9��ZW������}�>��q�@p��ZE�e[i�T9��L�1,���r����r�״_�u��v/���p��>%���XړV�W��k�z�w��o�fΌO�ԁn>�0�싢2-I��-�w�~�zm@o��#�Х�	��Q��fk�WW93�1�����סQ	�3]�-=7I��]'�͟RҖf�
������ �LR�%�7@fQ�;!�aC�=���H�Z������$7ނ�B���}%�P>�Ѳ��8]C\L*@�j�0@2���V2}B��<�TWCjx����t
\�2��I����Xy��,�.>��S����HYч�q�YT1v��O���*M��t����_���D��=���_�QP������)�滘�h#���%�{�oГԙ�AS�1^Y���!y��"� �}����q.��)�E���?Y��k����B�Q7�M�r[����=	�0!�8;���:Z!��h�g��>����h��hz;!R���0���B#�|68�|EG0���{t(އR<Z��3{�N^��M�ٌl�Z3$Ae�!:�e��m�D�?&�h'��,
���F�W��bx�l^�e%uSC�n�I/m[��x�V�R�'�$�雵�܆$��hwjY_ٔ��qC�xtYOD�&��R 4�� (i��ե�!c��/��uV[�� gF��7;Z�V��b�y�kG�pc
1,�2��{��"��M"���zu��n�|��|3�����QOʯf�e�e�����Z�ޝ�,J hy��9��"@	L*9ej9�:�����Bd���⹏:���0���Bf	�V�T@�������/Z��b�O�r��HkCEuLѡ����_��~�36=c,"0�����oG����?Zw�.�w$P�{��ڲ�i�lZ#�������`h��C�>�q9�VD/�B.#t��(�$7�����	��`��@�*�-���-O����q[�֕)����|��eUr�9R�S'�Mu�~|ts����5Ȯ���X�%J����݅�d�3濋�k53��.s��8Ey5�L�FT���];��K���9���5A)E����n���X*_�}"�@�Pg��:a�vSw�dQ1V�i�ƵA6��
��7@R!�)�Bm��^X>�q�x�I�]5�>qM;�<(`�o"�ҵ�zK0J�s&��z"M� E?a�s�"X�ۥ�R��k0՜@���J�I����u)��o(�m]F]ԙ��3���&>P<A�S�����{L�ӎ�;
���e�JaVt��O>���B(r��]�X�D�v8�0S�G��H�m L��~��P��Ea�G.���RPh�hln������p;+�<J��#��z��Ec�8��r��@!E��ݾ����in�בIx'����M�(�%���"�p���(dK�a�`�f-70�%�;�ˊc��9�7.����Wƙ� ξ��|� ���2*��e�.NԬh *��T;�
z
r��~�CCE�S���M7E"Z�@٭�p�Q�e�"�'�`�xyd�A�#����>\�h���� TZ�l	��/whf�/��*%�G��<�Laa�q��|�sl�sN��/���>�I�-*svRY:V0 ��W�5�}�A`C�r���96Bۡ���Z���Ċ(o�����ڏ�HuX'a���"]�LJ��9?��'�=�o���w����SM?�B�dR_�vo4:�������_/�<�i��U�1�¢�y�?D���Z'}�o�-����@����������1��ң8��� ���s��ׄ,f��1=�n����v� �B�d�
SF�T��c����L����S0&�?kA&��z"�:��O R��YD���y��[�A�&cEY���0٘4>�>���DJ���W�%�]�璱���>�C�P�����s�!`Fi�b�&f��2Qֹ1���(�]tu�9�Ju�q�Z
�9�]T9��VQ�Dj�Q�������$���K������QN$�+�'��(���S'6��i��Ȑ�ȽdP�POy�;��΍=�d�v���߶n��E����Q�R�$9�n{n(X���Sk%��N�ߪ5)�3�(�1h�������}R��1�㤰�8������. -0r��q�������K(LC�?Ki��逫�t\ɉ���u~�oFX"ؠ5�ς�Ls�#e}����l��V[���<��=���Ǆ��{Ns՟�D�0A )���:�'4��~��vP�ޓm�zi#�rhȃ��.�u����ެԒ3��F�����P�v�؎��r��Q�{�E�l�KAo�����AO���������iQ,/�c�
�?��F ���>�F�'m�E�ƧN��頍J \&̕�>�����[HD�A~�R����R�N���O'1��P}|'� �+�W=��2:�����0��	x
����L+6�H~��T�3��\���9�OD�	��5���_SA�r���3���(YP5�( ~89�U�V(&]��~-p|d\�'헮[��	m�)�j���@��~�J�Q�߭Rb�)�&B�z�X�����������!me�6����(��	hɠ��k%�8Q���F�Y�aD�0 ��s���0�N�cI�����&@���8���}1F��t�U�L�C�?/��?�נ��Ͻa�Cq5����J��}L�;Q�q�<�_}�wFcj�c���{\�̄����u���qz�h)��f�M���9@6e�;r�Iu1���A�ۧ�}n t%pfjԏݞ<��9�.��;H�w�YшR�.�{�6j:�1�b��g�$�H�:��=���A];���%f�`�EQѹڼ����Gn5����]�?:+�Zl=|�LhۗU��9�|�ȧځ�_�JQ$.{��R�\u��!Zu�z��P��F��L�*Z�tt@�6�ɐ"��}"�ٚ4G\㣵	>*��3��>5��:�8-�4�a
g�/�`�K�؜�M��~�D���������t�vQ�vJ�o���D<���M��X&��Q���b�2|4-��Z���
~�+`��;6t��]�
!Q���ع�����^q3�S�0��a^y؏��\G��a�������V��D�8�BIrA����IcOL��8K5�;����m�} �#�L��;(���:���;�Z#���<�
�V6���c���zZvoC[W�xZ�p�4�g"��,��\��J)�Σ�������I��|�N8�R�� �����G`���Qv�Q�����{��5�A�Jr������"�fS��J�4�h�S�bZ,��Ft���sp]�Ѩ7�3�A4uQ	��,d��u�l#͘��.y�/��Ĉ:��ά.Я�m\o1E��z��7�l�@߫�lk�Y�z$����q��j6���̾���ql,'�Bx�_���=RQ�䰕�
�T�D��-9Y���������Zdȩv�{fscL�Ӝ�V��ӑa��x�s��D�1�9P:��7efc�b�g)�~�.ݱY�����E��+<���ѝ���W*\$�m��N��t$��,��kĿ�ڽM�Ac�˩�H������_7c3�6/ĸe��Gi��{e7uƃ�IU�S	�b�dB���Κ��5Oiɑ��m�Ŗ9����r�\I�Rր~w<)' 6s��mSҼh:fm���!�(��������#"�`�p'�&/�~2������?�D�7�`Q�=S��v6��] �� le%Ė&$t�6H3��pEN��|I�.�e2ⳑV�qOd�K��l� ���׳3)��i���>[��ip��k�~����]� u]���`����T:v�G�A{k�����,C�Kϥ/U��&�r��	2�3�n�{�X���ꔨ��c�YM�����prǮ�0��7;U8�%�����|���qX��|�Ǣ��(�Ղk�Oh�UU2l0JI4�Z��/J�K�j��D�My �ٽ"�����,]�p�d�h%��o�O�*}�2��S�O�8�~�@�Y��{�5���2}�������D\&�Ym�cL�v�h�a�'5'ms;�ǩv#�A3%ɺ.����0SR�1����Y�����R�������q	M��	�3� �a��ͅ���#�߄��o��ec ��+��o�{9���م����o�|�S��|�A�&m��O>��E�r�~���Z-Z��--��P�ś��*���c�o��/�l"$�j2�m& ��H��Uj樲=Fu�%��P�!,^��|cナ�	m�%��W�
�����V�j���]�	QM��©V�w��);�J��#\1�>DP��x���`���˲T7�~mR�!�#|&�[��+6��j�<}Kx���Ղ��S�b����H�w��p�6��Ny m�>A
`�3����܌��D�|q�1��d���W*cxi2y��b�^>�FI�*?�D
�`���ǳ�]��L�u�2	�"�0��ݶ�I�_.�G�Ae�`N��޲]�]NM���|cD&^6P�F�*:Xha�L�]��_�'�ۄ�y�u*�Q���N�R�{Gq��m��?��2x���G�����f?SM.�`�T�*E�oH#��TA�Q�!q�r�!���P��@&�R^��~�M�(�����NK=�.�]��@�
ؿ�4�c@lT%vf���A�ݍ͹×�+�o����,"�$_:�J�׆��*��e�a<����tg��B�* ������]��P����}$ʙ���%���� ����%��V)P��l��ra.�L4����};��|�۩a��l))��VZ.0ӕ/�O�(x)V*���V�mF[�Z	���L�@) s�M�c��ټ��{�k��i~����bDo��b��%���S!�����_$ݨ���Yg�۠�L������kYK��+�x�4bv�������ˎU<
V��8�[�j��{/JҨ�����x"0n�2�������Y���Z�W/�dU3��������%��_���22�G�y#�BI�^��,w�
G�YL�j���bG�i�
cm�4���'���<�̩��i��c�^�Ǧ&��.��<Rw�1I"#�9�x�Z��F�[N�
UI1e(˱�R�t����g�����7m������-4�dvω��h6��9��Y �O_rP�l)PWP_��\���#L�ѧ����W��Hu-dMPR%��=�{KD=|#�?g7p��{8�or�r�;pLT�*:�k��H���� 3J�
������V d�������=�m�}t:XǛ�;�����8��}���F�|ܷ�<��v�h}��1V'kO]�
	 Ꙩ�S�8I�]���PG�:q���.D����0�*�𭭱�X���S�y�Ru���帱)�hV�J���뼈�_���}���$k�WƷCH�A�u=�Q�ھ�����r�Y���T�b-��N��E�0�^��򃥸{�W�4�U�8G�
���"9a�FAڶ���r��m$Q<(S{R�t'ևs�3 �
m���j�>�>��	�?�84��è;c�E�N�� \<S��s�UӖo]i�`�B#yG�i�����X���l��Ӑ ��$���>i��o`�3Ą�y������i�J�p�a\�ؗ��y�5�&0m��[ 
�a=��d����Lc�~�%Z�ޮ���M�_�-�8�V�W���y�N���k��j$�u�6����������1�U4�9��A�
bK!a	P��	R<&/���J�����(hwi���0w1��2�Su�y���P-� @`�
�~�/�Y�q�1c� B�l7�y�B{�"�����dנ��
|�ÿ-���6:�H\m^�Q�*�w9�3���<p�2"��c*�KM�0!�:��]���y���=�k9��z���"�N�5�n�/Q��/�Lu�/�ռcjE�Lꋘ���BK��`�@;߬�קJ�4d��7�>�|3�Wz��K��� ��_~7O�#�S��m���?����cB��a�
џr~��m�9������H��~���Ŕ$��WͿ΂�0_b��t8�����>
���d�z�h����pK�B���>����t�n�T�3A|������� �*��
��;G�o�t�ޚ����)���v�1o@���jGV��#J-r��6����0#�`z9�y����)���\�'32p}i kk)��\�<?�-�;������77J�C�pRw�*�eo&G�TN�����(�{>�ꖘ���DD��	]�h4���lEA2!!���5���P��^q���/c6��c?�'����3�{�������c�6rgvT>��E�{�\�y���(�xj�Tc0�P�l: K$x�!�J,H���>�;X������-@��e:�
j?��l-]����G�x9Z~7�@"��kEpg.�Y���Ḻ��Ir�/[�X%����	��wÙt>E�ο�i���D�B��k�&�|��D��o�{����&&�{�}���K
J�&7Q�*"a��1�.
s4��׸f�2��B��b������4��ʓ;� Sd؉��r�d��q����?�D�j��Ѫ���E�$s&|ˑM�E/t�.����(�nGP+�
?������;k�)��b�۝<����L��ٗ bWY
u[nm��aU
#H��G^��� ��F���A+����5��W��@>��4ҿG�W�����Ŭ�l�zR=�yf�rgi�s���JMW��(a�����LY���e}ͫ��_;��dS�`��A#CC}Q��c2����9S7X��Ъ��ˣA���^	 �VB��%�B/��%kI��I~��N��0�A�ƈL�g�Q��Qu����xY�.����&��5�I}�d���q/��y'�Y�90p����%�;�$�"��҅Un��_R�=�j�����z����兲f�Ud�J��9z���Y���_ŗ�ؤ��i�\����B������e�_D�@�DTyo�D���{�+�@���;X����Qr6��Ԕm?��������R����l��-��'��vrD�uo����� 1�a��cc)R�i�G��&WzV�]��ΐF�
eZH������ܑy�Z���ʾ�1=��D�y:�@6:����G��X7s�_d�г8�Q�r@�AT7�>R���A������KR�2������}���%�cA��_5�BiML�Y+D�C�	*��F����>�<ڸJ+(:�F�3ĺ��	HT(Xn�D�M�ı#���Lս6�����Xh�dv���D���]�s�������k��E�@Ux$ʊ�<��+Y�V��3��pF��-������Z ��e[c2!j2H���?����ɒ�E%L��	K~�U�?�LLr�I{I�3[=�e���j����n�\t�?��)W�2r��Q2c���Yf�����CY�͹��`��Ŷn��J-z�f'>��*������O$ǃ=t}�����׿���;&-3� ��,�m0����W"�T��*ϫ�v�a����B�y,�`۲Cܑ8��M��zrf��i��(F��d�?�p�!�o4�|��*6g�ޯ8���'�6��ࢸ��pɏ��)��;������fX�a?�b#�� �)�[�'�OѴ`���]�1=u�"T�z�z�ܘ����A[��� C�\�F�*���xS��Y��5�Y�#��l�&�����>ʑ>Z�.MX�g�|��Q�8����35���^� (0&_���� z��V=ڈ����9d�x���j�}BT2��������Nq�砑�u��a� V���:��_�df��T�!cO�d�m-��+�h�h# ���n�\�6��7��/V)@�3��:H���C+!bF96;uC�r���9u/�s��J����°b$�̳��/̏�o>�% �Γ.pa�ϯ�5>^������s5I�Y&3A�V��,&�1���y�V��'�:+2��ص��d��bɑ������BH�ZK���[C���!�-��,�����&3X�}���E�����|rK�+�7!O9��^A�TeK%�-��dj��`/u��L)�ę����=D���o{�ޱ���5�8���%�=M�룓���lK�m&'gw#���a�~��)*��f)׃1�z�,����S�J0.� ]A��O�FuW���n8�q�i�����.��Jon�G6�wf�a��A �u}O|	@��}YS�W�>���!�Pq�7�R���M�����o�b�B��ۂ��Ըd�~�p$V�l�Z�*��1VR;y�rT�f�(�@����r�1!��-�u�CKϞI#�M��H��#89].܈��>�)�J���f?��ta�d�G,�gQ̴�����
�����%�)}
�eK9{�}��ߥ�4.����
�(2.!ۣ.��i����8$-�>o�f ��H<Z�EH�~�j���)͒{R�K#�S�0D��Y�a�N;T�����N�o��bPI�k�|�!>��x�X�<=�Һ���x�(H+x.��F��+�<���!�BQ5�lVUn[�m��9� �J��TL�G�&!��{��y8��͆	tg!*k���cP����'��驸)o�;�ƴ��`�I����?St�30������J�Jk���)��]^vbm�zlJ���սF ��:mSй�w8R�vWf'ҢH��q� �!� z�L�"��X� ��@�	�3��G��s��k�x��ySo�E�a�L靉��Q��x)�@Ӧ5%fȰ00��]3�,|��&v��tZa��Tvuʣx*zA�K��o3���*?lN�HI�`y�NN������F7��'��#��	x)a���C��[�R<-7H�����~��!�z�Ar� hV5u?�+���df�w`��>�w~(����ު2�nk��W�����H�����Tt�P�al� ���s��iT�^U޼����M�<	p<~`�֛����>�ȪW/�[71��C;D���X#�����(�~rDE�M��0�p/�����a�'=S�\~G.�VY�j:�|a/�8�A��0'D&W0V�a�t�KY��-O�N1���9�������E���^�X����c�ǃ��V�N��@n n�t�Q�X�q[y���g��o��zxׄ���*}m�l���>���E���X��>��=��L�53#��5�р����Vu�IW1���c��̢����p�5w�w�INSfz4Ӱ������JS=8p�O��V .��M9W�j[��r����/A�A�K��S����[A�;�O1�[�ą.�����1�ol�<�s�*�nsF��͘~���wznfÝ�"t�ܛ�����[���~,�iwp�Z1��4f��b�zz�a{����CC���JF�{���i�7� �F�R�T��4s�b��vm+�,[4��b"DN^@�PP�wJ��A��cэ��yz�}�
�a���%�X����Kl�l~�+;�%3�@�H�������5��W���ȃ���P-����|����V)ǹv�#[[���/������D�mŜ8	O�~W1�(B ��:EAlԑd��@H�}-�9	`�s�9b@�t�B=쥽z��z{!3�r܆ي�K᧵$	������b�"��B �>�xsj��A�ko��?y]Q�%�v�Y�Q���]�͍�5��e�NC��5��^RP���aFq.4{�M�����u� ehz�v<LB���y��|5'�C�:c��d0;��h�~�y*�7����r)�yH;��4�|��S�q+_�y��4�{񙔻�H� |����4C!�^����N�;��߮�����
܃��픁c\�Ej�=.���f���n:��������!.{��G��؏1�d�y�Zǆ���K�D4��2�Ady����{�O�_l���)-8��y��x���v1��,�4��a�D�Z
�%�DG&px��|c�
Yy$�%n��Ѷ ��	+�TQ/3=#ɟbm	]<ow���f{�'��~,�̉��N?� �Kɶ��u���n'���Ȯ�	�G<���x� h�B�	�����C�I��w2��j��G;�ԅ����~5���֭�����k-�~qL|L0�o\�7��B�2l�Y���I i���w�ۇ�!�2F�M�a[��V":��B��L�T-a�փC����N��O���;F����n]�b��2@�⟥�I'{?&��II-~�pUI���v�4!ɣ��#Y�&��_����]�a�CaΨN+�D2���V�Ȯ@����Z-{���WdHH$!�<bt_��6\tT��>�Zw��H2�:����ā��
�5}�%_�X*:��&��T�Z�^x����OO&-�g'3!p��[�?��~}�=N,	����@ñ�����;�c+C��M$�pn*�d�>�]Ǔ�J���g8�"pȋ�����4����F���7�D$߳���b7�J����D�y�]{t��(V�$��+�9���;��-��!=���3,�rg��tDP��fB!��<݃�0S����U���������2�����,C�ϯܩ����4�y�^��J���F��¿{�<�
}Cn(���_Ec�IF-{&�w��] �2�х�9gƅ�u�`.�@wYFtIA~���V�+��y��4Po��팦����zR��P��i�ȱ<�e���AmT:5]~X��;K�v3�?�X����}����3t&�@�o�૬��/�	�h�՞ZDA��<U&^ȕ���}Y�H*� F���x	p�RJ뇠VǳSES<I)lL��1�;K���A��5M�=^�,����,9G���E^��@�/_��i]êa�p�U��2s��\Я�('�})м��h�9(�'�}sɔ�u��p+�qX]��QU+��yg�of%��7��cn�`;�yFDd1��f±��W����a+$�;]��W�P�o�[�<��"��*�C8A��R߬	�<[�)��9Ze��U[���B���d�o4S��VH�����O���Up�\ׇ�Z��e�XP����7)!%���;l�|j�؋rN�[��х������N�N�����P#���g���)�r�P��E��(�رY�im�ӧ�_Au�82�����RN b��h���
���ѹ��M�N�G�'ں�y��O�>Rm��X��N�̦���G��C��J�2�$��N=G��8��x����-ی�� <h���t,N�؇/6x��B
����������ŀ�H�W�jv����%<���o_���1q����ϊ���R'O���S����Ԇ;�=d������p�c	*Nb!p�1���
(��h(��T�������2�����o+ӂ�9=vf�6�~� Ư���~U����U�z�� �Q/!�9D����3��p�nB��$ȓ'CE��Gt��)
]BRYa�����mʗ�`G_a�x� �{^�f���x�6��,�,�d]�f�<��3y��=������k��3�m��]�x�vAW�3��Yi��9�H �E�-r*{���v���S�Q�;:��**�[�R��V��I�0�?^�m���hB����G�ԥ�䣃q闱���X�<��\����뇦FdbY4y�l��u�YX��\Gxfy���2Syu�G�Q�F�'�[��y��ja�qB�4��C�(f,<� '!�I�?���c����À�s�z�����J�cr�>2!�P�d[���|���UhfL��l�hzM�1)���u.$ :�&�`����UA�\u	^�x
�QA�&G�����ǳʃ.�5��x�`�SX��[��Ų&5�,ё^�Tj�ܥ�jO�.�T
 ��`�xܸ�����O X."v ��ՀU����.���)�S�~�)SWf�5
4Macp���S��6�PF�x�7�+A	C=cT��Ek��h��a.Ȩ��y�U���a���r)p�A��p�~�[�JM2^�@�B̽c\��;�XJY�jAi4�P�yTm����p�[��QU�49;/�k�`����n���!4%HS���*m������������J�ؤ^p��Bi�Gb��-����c�S�����ao�eH��(R��`~c'{:��� ���Ij6R�>[�������9{��5}��91��
� �$uֿ���AL��k�U�_������g�j�=�)����TV������r%?��IX-Blˊ�~�)jA�
�A0F�:����݂�D��]٣m�D��;&h������}7��X�ݬp� �X����N���������FH)ٗW*iw��m��w�h:�����C� j��a�\o:�.-pJ5j^u[͢�\Y��M�I��|<d�mK������M�&������#{B7��G2>�dI��k�"�
�X�G ���G[(�$MD��O׌^Q6�)j��gN�FQ�L�e=U��Ğ�at�S��2���v�\w�,��yB�/]	�x[�K����e�`��џ"���="@o�����{�yKH��KJt�˫˩����qIR���fB́krJy�#ꢄ$�����R��R2{쏽Q�}�SGi_�5�	$3��x�x�F9��
��c�H
WiUT�}�y�@ir0zGE?m.8����'�!���ȫ�|���>���+$顯H�3���Z�o��Dx���mV�[z�MN��{�v��!%���-��E;qm^@$�W�}D/����dp���3Gm�W��FF؟YF/���PL��j��h	�n�&Ţ:������jS�C/�Ѿ;���'�:>�w7y+t���2U6(�#f|�phtBg0��|�X��J:�]�'3/z:8�����3�E�8��j'?-����8
�L���!�yY?�ڗt�/4�7����սr�OɿP�GЉ�*�U�H�<�h��N��7=>��
;���7��@��hm�^�Jb��Z�� �C �d�B�����p��Y���#3��*M�D��d��eF���&��P�������'0�-f�8�H�>|dc&��=,��!k�ƕ�����q����~�2�0�	N�>N���ҝ���<f� ��j}�4&�yVT�F���\�'���D�N��7��0�!��脃A�Vc��I�J>D#*��@�h��BH���%Ê"#q�eل��4!��S-m!<p��x�;I��D�\���})��s���e]�*kw��8A�sA�+�W���ez@�S[1�Z��l�yYp�Y���!�&5��k뇒�9L&�ҨX'b��H�V_�]$:�����m �ʅAk��_����m1����"0���������p��$-pB�B�N��'�l�xJ�B�/��o�=��a(�����tZ�j���<�+���9`���\c�8!�h�;GIG��'q��%VXyH��䲡�L�Q���O�7s�2�w#��LN�6�hש���}�o|he￿�g��a�0��c"��@�o��r��N���Un9�#�{��
��2�/��z�������\�d|��"ܠ.��nJ�o�Q��]����9O뺡���`h�f��J��[�Eb����;�`3+(yؽ�ո}>��e�9z&蓯����A0�Lg$�Wߌ�	�,mڌ�[�p{���͒�1�(_�WB�N�D����+����p�����c�jWɝƈ������ϠL�9S���S���0�D"��%��f��/�&�e,k�T�v��q	w�7�?�A�:b�#�S]������Q�'���[�h��̮�Ǿ�kWִV�،+�Z�%�E��ֿr;��B�vY���n�b��;|�h�8
�L,	h�V�2���9y��x�n���$xo�Mfw_���ARl�����0̴�ygmm�h4�g�' ʷ�+���y��0��]W�V�밣��	V C����J�T��*�U�_�Ql{0B�KL�J*���R��t\�|����?Fӂ�����y.j"v�-fc��Il��_^�
�Otq32Di�7����t�����O��'�u2;����� �[BsR;�u5�}Y�󶷁n�<X��´ZƖ2�ܚ�Uc>׳xC�l[�i���e9��z�mۖ��*�( �/V1~�ˁ��(j!�G�{�F"�1���x�4���fAy�[_%{��W�5mޮ����ݹ��j���m����~����8rNe��K�8�޺ǳ u�?�ftE��ȫ�e� �ߩ��>�
���:��4�Qy�dƢ�o��H�Ő��=�%aE/�;����T�g(�<���^�kJ�ܞ)���I�8�T����Sj�����`�a�x!A�tl�($�Q�G^�����b��LK��̲h�O];5�3e��qb��+JS.�K_~�&4=<�c1�Y��RVn�EH ����S�ț�mȬGVx�I��i�1�K�DJòǿ�ˊr����[��#�[fWT/B8&��ϣ�:{���G	�uf�>��˖����Ni[��l�'@�L����Oj� ��Х8�tϱ�7^��w�{Ȁ�B��f�ҥM��Y��i{b��2ӊa�/�&F�5����5Z���{��8�/7�$�?Rf4]�� �|�n�]r
��0�H�A�z�å)�W4z��*I����H��]`�5K����'������Ș�*�?�[Vup�Ú[ŕK~�C<N��E1��22v�AJ+��9��pc�-}:��\i�o��w��2n�c��f�{�	-�&+ܷ�?��&�ٕ���"\��(ǆ<P�xʨ������)d��?�Į����v���`b���Hur�c�p���Z���>��!�(�}��H3\�o�M��>j�n�l>�x��&����G�cIx�Sz��zC9�*xHw6*��.�*w�v�<0���}�k҅ VXQ>/��vd�N��.kF�q�C�8�2/V#�� !�r[����P42�QII	<�Ź�rf��ot&�ܨ��r�3��4o򰒮���yG��nb�E�����N*�$u��~�D�olO�{z�	[���y
�(>T�pY����j��ł&����#h��C��w�x�yp�d	H�z����������#�4C��:P���k�߲C��
��Lh#�5I���W2H�Ƭ�d�&;�Y>]A���ܥ���E�8�6s��.TҨ�οG�Ug���I_4-⓮XL��寷�Q8�7���ލ��O��a&���
Q��4��v�]?�-����9��wu!Y��j\i����T�u���FK�?���D�T�4���������0�2_���^��fI�ւ��Ғ���n���{�z���П"1�#SE�΂%�~������I���'|71���~�ɾ�!�dq۱J�� �A�䍎 	5Cآ��U�T��"�&��&����q7��:�@��d���ǟ�]uz�u����m��.}��9�xɉ�|�[��I����g�Ŵt��dH�F)'��t̗�j�����W��v<fw�m	Iz�E�����1h�N�.5�.���	�"v
`E�_��ʴu�9s5��+pD덼��D8CZ�t,G��B@:�M�,]n�нɮ�(�ў&�4�F(ta���J��Yt4�h���CV|�{@��n��:$����\�\1 �'���|"幣Y6��
�iՇ�N�'�w�� �%�y�ٴu^��p���R�)*�^�sOݑ 't�΂λ�.�Yʙ�RR���1�I�|��z�c���D�A�?yV�/��Jɗ.$&e���ڪB�Y\jtVU�j��N����z&ќ��j.ސ��o���B�F&�:���7s�7%X�6�,ZmI�����3r
�+�RK Iyjܕ-1�����U�'�ۥ��&��Ο��s�>�1nf5�R|�pP����;�df�"�N��1����J��X��9�be�c��̭@�g��zn��I/�#��y^IA�zb|ey�"�S�r�M[p�P���k�f�#>���=Lr2�n�\Y?�d��d)_�Nޮk�e��k��?���������3wGc0��������*��I�vZ�>��?Ę �`�l�,�z�!� �{/���5�_�����q�-�Z��g���XG���.�s&K�l�2�cqp�Ts�i{S�GQ�g�]����l���z��"��lF E=�-��4���c�ʎm��
�t5�|��3�@���6��̰�U�������ޒh�I�*bzQQU-dS԰L����^�Y������0d� ��@Ko�</�r3'ip=���`��(Z�}D���̳�� X�W����_��\w������>�x�d{Gvuwse����)L�:��̡w2�3X\�l��s��ɦl%|��(�K�^�cѼ=�6A�Y
!g�����L'd���y��*�89�W/�Ʀ3R.|b<��֚�>]���8��(����"�
���`���_3X
OP����.�?����D�Fu�]���!��^S�߱�1E� k���e�h��"�@؍����V�ڲ�����:��_8_�<�)1�W�X�?����"�1DxT�ubb�m��sTQ��dP����?���a�H_�y��6��=�)�r��F�O��_ε�3�|���4c�[i������D���6����I
�fܚ���.=���#B��*�ߘՏ��0�V�?�;�ʙ'妭#��H���;�A������v+F�N�ש�fy����(0�Ȱ�<���)�����]9:��_ɹ�Vy��i\nn����OR��b>5�{�G�����^���Z�����S~���D:����k�Z_���-F�<�(t��C3�1�,�p��B�v�H|��+�뱼9�9@	J`��loY�9N��6����)j�	nz\���?R�Y
�ߣe�~�j���֕Jd
��^aG�m�k ���x�tT\�1��.+O�[5���4��'L�B[���D7���EQ{TY��6�vs��z;g0��؊�!�sS<>&��#o2u�N��v.UO� ��bυ��n�똛cc=Ie 3.zՆ%Dw2����Zl��G~Ɖ$�� F{h�tw���Ba��
��?+���cݿe���2��*;�����ڞl�@�v�R�( �?P;u�,�O͑�M�~ߘi�,�P����!�YiS�f���T����zSZ�y5��Ǜ?�	������ʩw(-��ӪRF���]g���([���|ftM����M>懛�Dx�p$f��pw@��(8R�����̬pB9,������5�{�BR
��E�*O���^5Z��P��Y��S� ��5(�0܎3�_O����zA�����g�0}J:�x������vS�U��"��l�ZZ�զp	��}�hv�)1GŜ�\��X���>3��2u9�lra��j��|[Eo�����ɀ̸e(Ef⛊���r����b�\l{�LX�3����|N�Uk���Y��
��z��Э6U�gU�/�/L��?�)n��M�utiʎ�k��7�] 5	35��ӝ�I����+�*��0�g�����Z��ݏ�
���/c��p칅���؀�%l�@8��\<�QE��˩ʽ���^乕�,cBK��i.4�w���PL�ot�E$%�����ڶ��h��=�W��yO��qd��M<n��>��C��h2�q{��_1�ud	,Ӧ�X��ui�����{�_��n�����:�j��#tҊ �-&�^�ı�/k��<f=:ȑ�úY�y�>�q�AX�ܾ�#��&_����C�u�!�4�pA����x]����9�/�tvxh	�j=�9te�úl�GE��*��U��1��������q�R��괞�����̾7~�m�K���Lg_;����8VJuM��U��qB�s��@�`x�dܤ��G >�U溧x�q�3:��{wP{�����<߂H�/��:r2Mh?I��|!qF��'��U� (A�N�"�� J���;�D�K�1u�j�\
����J�g�'����Vu�>��2֨G@f��I���.f�Q�F�0��+>�k���ƃ:�i�䚗T���L!R\���Ɣ�F-��SF�C�=R=]����¤R�q]� 4�����R|�+������n�"�~�7�|��јM�"��=tPe^zQX�����^�Yۘ,ӝ���CM��Ư���*�Ki��Aq�4<�_K�
��˪���fa�M�N��n=b��'p��	��s�>Od ���"wj`]�p)�[�if�ӄ���ά�!/�Q����_o'r�N�y�����X
�4dRfI=vm���#��	O�TEp.��\
��<#�!K�U�ō�{g�U!`j'�*�JA�b��Y�҂ߝ�ju�.T�b����1�~ �5���AY�}�0�$j��`�d9���sOp�"��D���:��9��ȟCC�n>�w}�w�7����g�b|�~��ו��3RW�L�NQ�^I{4Ͷ����@�����?�4�H^��B{��Oܘ>9#ݭ$��y(��\�sqs�s���)<��g���jJ�l�`��y;�tǒ7�#[��s�2�jʵ4��h Ь|��ҧN��x�I�,sb^��*�o*���\���f��w)�/2�@��@΅�tGf�k]E��5]�`�����|go��MGA`%��[<7�CRq��_���Q[�Ŋ�ч�u/*�k��W�NR|9�A{jpi��򐡰+ނ[fu�I ��c-#2��H' G��g������yh��:�����4�53)�Ɔ9 �苪2������N_<2ۉ�����	��A-j�`�J����]�='i{�a�������'�y`e�F��֯h��0���`p�g�r(_�p�R�E��Z��]����2����[�� Mq�Xg�0�r$��ѫj�+�����;7�9]�p�a�◫����.<�|��W�?��7V"7�zf�+
6[�X��� !��,�h�pu�w+��,����J�>=V+Y��"ѫ(�SC[`��jM�,������)Wβ��݇E��p:u��X2�se���'t���w�$Q�tp֝B[э>7��2:�s�b�@!f�#��;�b�K0�m0�n#V��
�硶^~!�p ��i"��ܷ�n5:(N�M�^�\e!�[�nm���Q�'G�*J3�5J���淹�U� o�mYm����߈c����q�d��y�E��3����˪~.��>�$م�,}���L�~y�L�t�(����;ײ�&�[�H��̘�o��-r�t�D�QG{Od>w��rC $o��ܼYу�^�gP3r���e��������U�UrVUW��Dd1����kb'7��n�/rL��s�%��^��n$\���cŪ���p�Q~�g�����K�0�'^�ϔZ��;u�"�hq����V2�	�gM�:%1�U��f��թ��}�# ��3T�e���\(��<0d��0�l'Ϙ�S��|$�H����y��wC����n��#�#'&h��v�j���]�A��̒�>�e���w1 H�bT��c>Pa1��:"PV'T�-Ƚ�l���&�N����׺�g�OnO65h	zY��z�ۮ�b0�H��jc��G4Z�ۿ�7ZG��=jBJla�M�� _QL�͇����Y����4�P��QUc�8��_��[��,���݇х�w�W��*�[�t���'Bb�m8�y_�	�� �U�6�@����[���}fRLN����:@N�K��g������UF�����q� u{�Tp�kH�lp��,}���VÕ��%:U�8]���~ �Ϡ)�I�~z��0	�_�N䚇��a��z�K�y#��s_P�6L��L흭��u� ���\eDA�|,���[a�@��W��H�x�����&�IO�G�dk|�^���~3������I��A�"Vm�<�ų
�gQ<a������]fQn����
GIٷ(z�#����}�kClK�If�qM(]Sݡ�P�r�qq���dmyd�.�x'�~D(��i��*����W^���k� �%M|b���縤��{f�kjqe��l̤g�su7H�Q��~|ŏ���ѕi� ����JM|>A��w����U���1\��IsA*^a�����A�Mn�M�O牙~H�_�n���^.T%�Y�
���Wa�-����
�F��S%�n����YS�qB8	�Y&?B��k|[H��ʖI���+M�"\@�WM.I&�n�u*)�����E�9�~� �)v���Q�>"����=�X�d*?��5���+~���􍛥���[b3��Lb��$A����(r��A`�nc-�	8�����r��� �a�H�@*�D��n{�v�pJ��\����v���
�@S�X��G��dn!�7�y�=��By�{�;W&��b�CD������P�oYd!�o[��z��5+�y��R�zG�C*�E����c��s<}SYb~��i��}b���wt�L|��o�
"k��E�6�����
a�`)8�������j���]�����z)"\�{�b�F�s���A{���xq�L����"�9R�$��*����]h-N��&���/�;��� �h�ә��3+U������a��?�rI�O32-fG���L����2�X�ɯ�j !-;��^�q�l߼5��sPD%#Ol��ź@xf;{3n����w��UR��.i3���D�z�lhID�Q�hA4\s��1 ͕��yZ�]ʧ7�
�@�Yjub�k�x��*}�(��Ën���+w��A����ޛ �`�j��AE>�~鿙a�D��2��x�M��C3z�w����nh�$��n���	e��@�U������EQN��T�Z�G/Z���>�I�7�~�{��͔K��ħ�e�D!G	�;	�$�yn9n+���t+��`�lp6f��-���F 7�(�19��ܳ၇E��{~�_#�*�S-0J� �͛i7�G\��;�U����6���2T/�r5���mJ���
�iou����3N��{�����& �а�0��&N�����˔5L���[�B�xg!�hŭ���ls��m�G��� ���N�p��9Z%Y���?��*K1� ]d��ק{5
���ŉR��F��݁��n٫D���X3�]'� yo`S
I�p����@vK��렘�đ�7�F�7�^�I�'?&c�c2J���G%�1��,]m�N$g�p&���5ޥ�]cN> � �#���~��D
v��O���\/���Os��a����~���S6gX��Lt�ߙ����P<@���5�p(���2jw.��1�^��\�mdF|�0�s��2si�O�څ�٭�;9�r\��f��UQnP>dn�� Y�o 
�ަk;=�zM1�x gm�yO���nw���Ao���2Q+�������@κ;2Ga��'G�N��:�P�
/�e������?V��H�+|�Df@THZci*��P���;q���qY�HT��Ѿ:��}������+UС��$�7y��w�{��ݺ��+*�΢�v���6J�zx�cI�"��{o�:4G�ޝ�u+E#��Ǧ�s5�ZPD��O�;Ĳ��+��fC^+pv�m'�_&���һ>Y�3k�cp�R����Y+gؒ�����-fd(/����Б�!ap�b�� ��	{e|��������ѓ���/)T��r�����>EL�n��37P!�Sc^�ߎ&O�hV?ڵ?���ЇMu�_ǭ��ke�ۯ�F�	6Q%Ħ&8�a�̖� �"s&Ĵ��I\��2�qx�D�����]Y�ATOs[�ɇ��U�a��U��n�Lx��K]錏9�_�q@�X�v5o1�2��K�"��A[�� ݍBɟW��!��)�)D����ن_B�Y��'cH0_H�h�����ϓ8J��;ċ�}���B���S��~��:���3P[�����0�Ya���f�.�#o��)�˜~�}��I�������SE
G�K۶�#�u��B�ړ?�/)4����������p7Y�􎋉��\)?��[nB	Y4Vl����+D�d:�ԖPGL���;A"�nF����x�N�+q�wC`U��j����n_��2?�/r4э�̡���?�?<2�í��f��v5�(´��~w��>����{��F��)�V*w6�@� �����>�2������&vIo�C,�z�ጇ��7��Cc:��Py�:j�\�N��������C)��%�6YXD���Xs"� ��r�S���Z�,4v�uy-_���&��G��W���g�on�r�n�"Q��߀�I�1IP.�!��F���� �'�]����t;R����"�-%_.���U��C��q��W�ү�B�O#(�&B����ݬKU78>t�FM�!d��s� V�Q���D�_���=+�$~c�q��
����n\��s��Π2A����$��`�w�C��dD�^]T����Xe�u�Ra}��MI��Y0	N\�ru/zA=�B�#)vf��:��R���~�ۇ͏ܻ�IM4��E�T�|�j��Ym�c�
���>+I(P�ǀ�5ɝ�t�~�54A��╊��qF�N�j�6�� 6�g"�L�X�YA+�p���Zga-E�(g�1'
�W�E��դdo�F�g���l��nK�:RkQY��� 5>z�<(L�2#,��Z�)[
�"tF�%�h�JY���jz�zYgt�ᬃ�x�S�����Kw���Pg:p�d�ao��E��Q~@��K��) �3ؗD�� &&i��`>	�7�ei, �
y��p&�[h����R��ć�(���H�S~m��׸���ɗ6����AA8L/�<an䧸y�LJ�([Ļ��1�t}�"�P]�}�yX=mL,I���ȱϱ7u2f\�[��TM�31������$���v�0$ix�E�vt��&�S�uF�����.	zI6�;���2�m�@��n,� NjK��` � �sR�r�@	�\���+�A�|���z�5.��ߤ��va=)=0�5K*��G���Mj#��W{}���w�CV�ו�;��v�q�EK𘞩V꤃)]�̠�:eYF5ɥ��&�S�[��T&��س^���@��A-Y�a��5�T�{�6d=���Vz�Kl��S�N�S4^��ԛB�������]^�g�W�Eym���҂2�C^v��e�~'�P��8�o��?RDp��O����_H�M���3�}�S2S���#s�|}�i���p��r,P3�kud��2��@o���7�H@#�Y$P�7���G5@ !p��O���:O���T7�MY�N��s��.HZ�O���@:��f�hp���N��]�����b���~����A@m�k5(��g�?x�Z���)	V�2]��+��,M��Sco��CKI[-e��0I�l?WR��>���i�(xF�zf��h�����,m��G�7�����������Xg.�6��&��zX_�Ƒ��M��O�H�gh�p����hU���R���qU~���L������Y�Y��b�2�lt
9DO�qOW�%�f��qY~���N�A�۷ӂ�)���#	�������� �͌�n)1�޼��L�D��]�cNDi�'z���p�[�`:;i�#����K:�]����Wل{�0 ������5�c�L�[�.�41�d�7�%h�N�/�(x�ߪf�v5���5SG�Kj�ǰ ��$_��M��L�U�c��k�^�����Q���%/=!�ۋ��Zl��F��%9�]����jJt������H"����������F[H<�u7�d���K�Y)��c�q�X�j�i�9����0����mM��,\%�N�*�*g3�Ε�?k.��r���z��Ӈ�2�ƑO�u������K�c*⎋�b8���j���:�ˆ���7dA#�����1���V.��\J�(zj~'7�k�)��ښ�7p� �l*���FZ�C��D��ґ�;&���7&l�D'b8m
G(�l�O<����48����5�`o�k=��&�=0��	�Fh�:n����F�0|3q��.�c���-{Qކ�Q%c?�oM��I���'="����|bp��0C|�0¢���ҳW4ZϺY��7?&�' ��	Ň	��؆,�f������e��9���
�ؔr4c��h�����nt��п���]M��>��1L��3M+@F��N��֫h%�!s [��.l��ƾ�-O���=05�r��H��6�/~�p������[*����T��6��e=g�a�~')�S|�jq"Ä���q���<rٕ1�/�_�&x����`��I���R2�Q����#4־��������G��T��i(e.�F�p�9a�����W���,	J�;9C��+�U���A��E73��`��zg�{�4�C��R���||�M?M]��v�ZS�h�_cG���}5o�-���'����]{�M�!^	�032��v�s������ܟj	m�$�������6]Y���[���P#���2�G_�J���R6D3�a�p	塞��G���D��H^�.ӯ�3�A+0�$gX��gW���٬���(����PH��7t�%Z���\�ʟ{z��!йsTazE��n��� �#��z��m�U�>_{�&�-9c-tn����Տ{��C��+V��#�������"�Z�o �j2_�_��no�n��A��֫ƥ(����cHz����pX�&�	�?"Vm���W�6*:q���m��%O8A��U�5F6a�M$fy���d�B�_^�]�f���%�����-@egs1x1�T�r�GvN,E�I	g�N����1)��I����[��Tpu3�sJ:������V��W��4C��jb��K�F\������'c2�bcȿ�� U��+��lo����vh�>R��y�~
m}7+�,;�
Z��)R�rLQ|����0�2��w���ƣyQ��/�u~��$���s��x�<��U6�:�p�T�t'�|�bٖ��y�A�'��D��AV ��u�� s��ݓ�W��g�j
��f��aie����v�F��,�:�rm�5O��>ԟҪ�}y��a�4�76X���.�P�Y�F-z���;�|�JǮ�g�:
�ꔱ�����7���pfҫ'���l��^_X[0>l� ���P{R�W��݂��"���<�n�`�?$�%E���#ۨ� �~q�7��kWdSD�]Bwzw�1�Tm��c]q�ݶ�5���G'X��$��hj�r:���&��:K�:ƶ��p��jL�#�����R7>A}!�{��B���=�-�ّ)�,8������,m첇|�`�šL�,L0�9S{�Wi�G��gMT��π�թ�W銞�H�+;U��Adx���e�m*�ڟ:V}���*��X>&�A�W�ڿ��jO��:��-8˫I>-�z���qlR�d�:�u�٠r�s�^켽�UYNh�)MF�e�C�
�VȤ��s��$�k�3�cSC�A6z87���4�6l�22�ʩ�7�N��h��C���⓳�N�#���U	���+-���3�(�V)���h�����KpR5$�W� �61��j�����c�
��\��Vm��h���	�|�.�Ƭ��z�m��iSU2n���O��v��L��Lax�[��+�ѫ��vt�s����Icv�o�n!��G ̒�Mt�UUh(��~���jJ2�!��4�m�'v`2�>�(� ,@���Ct�۠�������w7��>nFN(�t����44'�ղ'���3�6�ѝx���=]2�C�2+/�m���4?ڲ8�Y4���d\Ԍ:W/�m�.Nf�y>�j�:��T#nnc:ߔ�w}���^߰n�Y�2"�'��yS�в�HI�F�e���6��×f(���We������1�A?���F/���-<�"t�:��B��'�Yδ��N��DvB��@�����:����7�eOMɥ�)%��,oL$��� !��t����U��'��!!��Sժ��W����An�nv �xy�Ҵt��Z�	2,��!�����tW�Ț�-���P�܌���M�-���!�U6z��p^K�k��|~-�` �(��9-ΰEw-"�i�6���Ҙ
���?P����%>�����2Z��[��3�3$���8C)�C��f|kjA�D�h@mԖ�>p�Į	n%2�oQ�Hԫl���(Y�ޖ�K~vy��e�j����4�!��m�L��) ���h�aLt@���2Վ���d,���
3W�J^�@Kԍt�>��^��9q0��ԫx������o"����S/_��&�>E.���͓XřS�e�-�8�w�H^�J<�n5 -�FF��-R;��po�e�a	jfDd�7|gi�uל�)�oFT����ަb-��?/ͦ;���T�͎b'���]�	B��z99�9OG�x��Y#�@�������-��[@5�dE ެ��׎��J����s�����X	�Mp�^�������8a�!?)�Lg���aV�=4��i��2��GdܨK=98���̸��ZۮA�9H�ta�f�U3Mm�b"�-���>+ѫ���7��.�=2m����ʩV�<��:��i����*�95L*�f����X ��ߌ�������5�2��p�T������!�@�[q4��� r���t �bh�:��	.ɟ
���&�/q6�^"��Ins^_?�R;��1?��gT[���N��� y���W�
1�1w����J�"Q�C/J�@:u�K@�C�2h�w�����~��8P�9]����u\N�� �發LX{l�Բ@�Y|g�vˁ��$��Ӹ�&�c�+���碌�U�0�B C�u�/���ϓ��k`8�Kx�lc5�0I�^�L���,����8M"l���xI���ǝk��{L~l�6�WH��nL�G��X�f�p��l�f����k��j�;���o��\M�S�e���%���`��/�.�T,q]� �d�i^����,A�v]E���[�,PJ"���WX��Y��m�L7�Q�fsJ�_0<�pq3��	�+��9Au9�C� �C��%F0Z�I����M@��I�J5W�D��5��IW�����q�@fq^D�Y�G����F��YɌ��*��N����8�����Q�p��^�&�L�:ήl��$w��|b��"�m�.`���֟����A[7��$k�P�̽*|��Ƙ[M��d��A%��7^��6J��k�X��O�8p^�[ 7�*�+2��K����s�4�����f��M� ����%Q�Si[��r�?�H��,S�9����F+Px�f���v%�U����m����rC��Ye��ZV�s��E�������i������3�K�����&iG�r�{��:�@�[�8n7�d�6g��(�Xi��$ܶ>��͝ĥ��J�gA�954T�/�����bm�w�ب���^�/�T�-�l�UEKk[��'���n$P�qCT3e�G
����׎�.�,���B2?su���覉��. p� ����"5��Bz�54���p<KJ���h�(�AZg-�x�	�}�-�MӜ�Q9���c��SKR�8P>�6�O���f�~�;1��{��q�� LB�;�����Ze�Ai�HcN[_�����n��lqi������1�>�!�Xj��yǷ 0�=��5�2[�磼��߼���:������{�Zr�BoR�u0�e�'l{�q���8�g�Y-�����g�!a\*lp�@�z��l!�k	��D���x�e=�����k�2���'g������Э�� �<Ձ�}�r�E��*w�����iӕ����&�܀�g�6��1���|�w5r�ݧ�ۅQt�d_P��2�g���=oyoy!��H���ц�kG�ɢ���[�ܟ0�7đpG�T�	kf.�G�͊�c��^�B���2z�U�2�� j�0�����z�h~&��!$5	�*��;F�lz�d��z��i�"kW�PMN�M�~���?*u��?���I)d�s�~�_h����bȭ�Bo�)�i���=������)�i����l0Qοj��UD��MR�{$�O��<.����O��D,�0���a��/��sdv�U0Ym�+oS�ě5=�z�
�����`dD�R�R�O��=�s��mȕ��a�֦����+��`V&��� ����!��nN�o�/�;���e�V��g-(i Ȯ},�(�����j��?_��^��m�|b8����]��A�� Zѽ�3s�f����,ޕ$�$BV��t�z�¾��LڼʇV���7�L7C�R�8&�$X���i�����h�GtԤ)(�蠢��l"t3�����҆R�I�7s���)>�E�	?�nټ\aC��R$�U��oQ3.����Pp�*f�D#�J]�]q;�rla���)h����-?׏Bx��kR�a�p?C:�̼�LژsYtYh���Ǧ��k��^v���o�9��u͍{<��	hz �,B����F�w:H�I!�8'3h2b*�I���|iB��a�L�pUaVB[Y|�7�D��G^X.A#�t�Nv�T�I���0�a��dA�Q�I���G�ZJ��
֫m ���g� �b!��h �T�;ۖ�n��:�ئ���s7�V�k�Ei�z[���~AU�n����#�q�vH�^���7 �##�Y��0i}��o�$�r��,N\�����ѫel4}5E%��g�U>I6�eB@w�':>n���^��FZ�C ��������BѰR������럳�[����
l���K���P�8��hH87��p0�޴U�-�W��R���#*�<�b�������U��:�{/ٕC�Hw\1���&�{��jC6M�%���/�1�PS�����<F�.�9p�÷�y#�+s?�* z�X���R�6�u�M���Jf��o�xRm��G��IX|Ec2���mނ?�s�"���oe8N$S r����C0u�e+�N�\ �xė�KJ�=b���7�����v ���k��'����ZĠ�d�L�
���&:#�n��b�ۗ�z
P�Ћ#��q"�j��ϱ�x�Gw��*y�jaς_�@�bz�0&ݜ6��sE)A�r��1�vX��ī�q�ە�ӆ-Bˊ-�ܣ���A>�Vri������-,��
<U}�K��4� b_wߦ�V�.��t��Ƃ���t��Ct�ل[J3,�t+��ު���o7�U,�9�)�Y�~x����l�;0��p��¢��I!��$���&���%!|��-�������۹Q��$�t�/[2-䗂��m#2x�Đ��P;��T�������� OQ꓾��i��󩙟��:���/���pHÅ�����)B+�T�&�{CA9-\�-3���_ ؜ɖ�p�Ʋ��g/y`'�;����P�#�4�A���!Q����D �	�dE����7�;
�,ҏj�=;����B�W.	��9����%��u	(��į6ܙ��<y­�;'s��gA��Q���oWo�w2�7.K�iZ�ji'_*���*x�8��3�Yl@#��y1g��zJ7X��7̭��Bq,�� ��!Vsm�#����J!�Y/�֘�v};詼�{(ڌL_����Ն���0���tp\�M��˿m�J���B5�찱C�7�?��v�n��b<-k*v�"���r5Rk%�x�~d�D <��qu݇.�~3��a���%���\D��!�?�d;�yW��u�EyԮ�^{�E�L�xU�����W�D��su)��m���r�a7n�����R�E��
l��dҹ����"&%����N*=�*�R��P��H�o�C'��);�)
���C,�T<ϵ�ħl��E�1.&��mL�K|s*��^\�>��ב!�����p��|�FY���g<�}ES��$Ǡ�s]�Llb��T��;d�D�T�Qv���y�^��-��:�+�2ˉ9L&���GL1v��t�41�b�юs�X��Mx0����.����. ��:�W�U��ϽYrH��CeQ��ك�Y`͌2�^�4����m�J8oj�K��,4���XK���j��������K����!����4� l$#~�%f�X@x-4@^���.���(�-�B�BG��ΗkCk��a�(�44�q�O�������i�5:�.��(M���v-�|���lN������!�E��	{�_v3�i=$v�=��?̓y�%D��F�������>��i�(bT����"]����ЕN��gG���۹�:(��]{u{ˑ��x��FҔ�Z���^s�+!�á�W���"�Bn���'c�ތ��NF�_��g27�� BA���tW��x1�;�+����Os &��Q͢�a"���LTޙ��c�W.[!��q�,��]vЦ��3�R1��2�܏���w~T`�Zqavt�+��z(���\�!Ɨ�*��45��Ÿ{�g�-Ncx�&|�٣i�	9d��g�sO=߳���1��Ydk-" ��z�x���Eg�A0�"�����8���� �͘�6te"��@�3�]a�R6oo��Ҭa!f��]�N|�x�L�����r^!.&%n���W^��k���X>��A�e��Uo��av��d�m��3
#��6zU���Z��?T�-�x�gC����O_�t�Rwl+�Չ����'�`2�U�^���Q�݉�0��Q������r	m�'�������Pd9:� EV��^/�J�,����F(�@�����Ϡ�;,ĢK�ё�oIW���\��o���.�FC��������Ͼo��������I��ĝ[��  ����'�5�h��X��=���4?���nf"�!{v�!��K:���9�%�}����!�"��~���b�ٛq�4x��:���=]�B�*z �e)�I�)�_�o0x��w�,M^9��Za��:I�)7e����4�� �O��~it$ش�(���h�=�S�0G5�A.�$Y(5���\���3mϔAk[����L�M���^׈�gk�����z�����v�]�^p�X�[����;�_j\W4w1\�P����u��,�O�_�ȕ3k��9��VC	��?�u�e%�#��-21Ec:��`ġ3"[t��6��\�^"{3�o�H�J��y��҇��Y��u��9�df(r!Li��o,�`�n���w'�|٠}
�����׈��?QJ���n�(��,2�rǬ��W�y��vf�T�f�<s�㊱�CZ �$�!,��b���<��~m�F��Q��~ye�������fM���h�EЂ�f���i=�I�g���;�a2��� �o�͑tL��y��ʰ��˚+�֣�X�r���l�R���(���hjF����J;���p�vr����ؠi���2}�SNVF%՚�D^&k��j8�b�w�m@6���/�����9vWx��k�&S��s	1$]���êj�:�$ycJ�Qs�|�Ҟ��V�4V�`M��i\n��yj.��A�I�ys�y[C��C|��G�}����t-�~eF�7U�$���5<7�s��2u.laa�P-�c�]���[^�3��L�Gk��*�Β���m�yB6�'�/�-��`�;�<�P�,��2��Mn)xM�S�'kz_��Y�}&xM+��:�Mk~8��e��uܒ�5ͬ�䍩&A�	���U= J!�$�YQ��X����4��1k����ch@��a�ȕ�����N����Y����n@]:5�6��%�9Em�x��1��N�FW���L	 ��L���M�K��mF���@���fM��	���L����(�s�e.�JO(z���p�s�w,gq��t�C��t2����Gڻt���/٩�����{�`X1_�i��RH�j�3�	���S�����
@qd�a�y'��C(�}�C�\���G�&,V���D�k�YvZi�1�����K��v"��V���@�8I���/0g��c_�:�w���dnhʩ����k~KAR�3Y��S�Ǩ	�mփx�X
(M-+�2mȶ?<?ENv���Y��_*nD�}Z�9���ח�����#�B��*J�,��m�clK_��"x� &Iȣas���Ղ��a��PM:9@]!A��@.�}@���[���~B�Z3���/-��y�a��]���OJJ<U%����=�cS3��e|Z��S�,i� P�%�	�J���vw^��5h��� <a9෾��y�ʒ� ���'��	�u~�B�[FԄb�t��Rn&�rY��;��4Gޚ�3�?����T0'�)t%�,־|\ۯ�����?�����j���}*`� jŉ_��sR��m7��E�x� ��G�j��RL�vg&�K"
�{yQ;kfh���=Q����t�u��Da�ې�G�_��S�xаϮ�Z�<T<6=%�7v0���!(ҀQ!�=w�<���KoQQ��^�n�*�%`K��|�?�@�;��i2b�RtT�8�'��(���zI$k���)��I�\vUe��=�s
�G���c�)���q	*��B�c��k����ʁ���$�`#�)*��G&?e���qa��a9�^h�2ȌAbO���ϵ��*��j����䩏� �FK���3�8ï(�xNd��<#$�)���3����h�rK-����H�y)K}�m�WY���؋P�P���(% ��|�ܵ��s��/��Mݦ�ǥ�df����=(�X��M������wg���L�^j�T��f����Ð��qm<�o��a���j<3.��w�\�u�0)�F��n��s8N�]%���~�l�j�j�̭=bo ������2�*��9e���$q.����B��r¸*�d��;3�EG���,�䈼�)�)m#�︡%�t�v��!Q�j���o9�I�ɋ
N��S�9�������M6)�P�.WYd�vH���BM5NS����D����H��3��'�3ǏNP[�d���l���I?�U��q�E�x��X'A
D{�����=Z]�T����u6�ժVߌ���C��*d�Uk�:22`/f��?�r�.á���~%�&n��˩�������L|���c�-���u#`�1�Je�3�:�YǾ�>��h�Y�3*Kw��G'���=�ϪC ���T��\��wE	/nk:�0��X�G�Z���,O��#��n�
5�@���5Sa�d8������(��C '�AL��+����]"�*O�g#|��ڤ�/(k؇q��i�e"�q�Zi��-A�H�c��y%>��-���D�->����zv�����ƻ'Z<ӭe����yQP6�@��d���bb1L�W!�w�xT���63�(��fq*���N<`5
5Nč�r_ ����k�ae;'���u��%�b��I�%��z�cVA�Ebi_�E�ؒB2$p����h���%��S�h������.{e�0�l�
�ҪA������|���O�b��y��`H�.{���B�X] #���-ܗK�g�Ǝ��Ds�ۣgx��Fe�+7*9*�?w��I@��F�Z� }�&9�/m���,]���M+
.�Y솯�z׫]��s���GF���Vt����c�I%�-�4%A��r�u�y�"��r�k4���`7P�&E�R�r���Y�ל��S�8�,�Ƕ�NmE��ށ�>?�ang&�)���;���C�+W�~��/b�;���eK�n� o��^��_�#�o�@�ކ�e��_��!�Ӫ�R�βB�>&ݼ���Rͩ�e~�J�XTz��i�_�=SaE!�\�c�qA?_�����V�r�%��R6�9�2	�cEs.��7=�0�WQ��r��jNX����7}!�3�}XrȞ��`GF�U��~x����Ӛ�{2ӓ�]�={�_���g��[7�(oP��] U�(W��o��no����W��IV��x����4&������|L�����=Q54Н�1|�
������`�a*DʱwOH��Q���>���#��M�fD��D�?0���b�bZ)Xƪ�.h����t~�5���W<���t��Z�&l�$tOZ\n�4���߲hpD�=ǦL��$ѢP�݉4��sW�Yu{,�dWO(�7�P��0�����_6'��k�)�H<�=�iq�~�u�Y���J�a��u�k��[B ��+8Ucppc����k�&���;�rډ\O�����9���G��m�$]a��;K}���m�#E��t-5��_�e��f w"8X٣��aw���M��
�7MLFi�0�sON���ނ���
gݲ�	��o��ϙ$>��,�5�FH�� >�;˩.��H$�{�x6?�h��7�ҶP�(�1��(S�%�Y�خ�F ;{4��Xai��eR:tD�﫞�1�x����	�v�d��B�4cq:@���i���8��i�C��. ���fͳU�U3��Ɠ�e��ד�	i6�S��ϸ�����He��8�t���[�5<�c��s�k�F ���r[O�N<�ʒT0�����;�L�$b7��
e�V<����Ue�s�ޕ�X��Cf|��,����Y%-�0)W�=��C�����H�y��oJ5�����r��Exp��3�\F�n��Щ�3@z"/�,x:E���D���H�
�ޟ������U��%n0��
���X����g�g��޷��l�k��-���/���|�~n����A���7<F0WU������IQt3__������=�iE���I����_���:^��i8��D� >���X�%�Z�63�de��l�v��	�w����ƕ�<�V���8�؇��f�A�U�7cQ@��Yތ�L˛��o�2¢��1�g�w�$M��i��HNq��gZ?gM!�$�ѝw`�J�7�t��B�ͷ+��L�d>X�_U�mtB�vE�Q4[<|�
#�/5p�k�8p٪ڊ�̱)Óc!�j՟�t�ݓ���
���g�0�h�{�U ��"'�����pEZ�P��C�#�������"W���f�VF;b�gǂ��\vN$�� �Ҭ��e��c���+є-3�WW�8�|���1���S�`S%�8
�a��|Ϥ�BfM�p^9�3D�%VAga��Y��p��oK��]��i�>�X��p��5r����T0�LM��]�ӷ�<0�����n�R��d���:����ݒ�:�c�/�u$�v�{���Y*���L8����I�vb�h6(�2g�W[�u������X��@�߹�-�|q��PS�ߜqon�	�#+�
 n6�c���W-T\pgˊ�fh���/s�W�Mŕ��%J� �-��g8��YZ�lP(�L��ַ��_w�`�/ld?�_e����*�o���$F��<���\2;�ޔ�8U�op|��R9ǡ��� ��6��n�᳦��I:���r<�ׯ�"�(�t���}��O���d�/��Xy�(6q�ά;�&ozי�+ڽ�-j[����{:�#gQ�2��hW�S�J��Gl�1�m�,���t�=��z߇��ܧ�F�����d���$C�-;�O �{�� ��%@�S�Fй�z'�t�c��4Յ�	�PA�j��f�Ǉ���^c�
H����+�(sAnz�z�Dl�Gk:ʨ:���n��.��G�%��hSU:�衿��&̖\�:��4 �,��&1��jV,�w0
([r$#X����$*tEvi�L�A},յ�rʤ=��#��R$�|�xu�*ӯ�¨�ꉧK����-�u"�f3Yp��
l!݃6��.��ߗ��/��u*��;��ֱ#a����7�^:��ȣ����g��+�ݳK�nb0�H����( z�޼�Z%���MY�XH��ӥQM�	I��/��B�O�#{wn�6H�E����K�W&������[�0�,��~@a}0�b���RC)
IXC�ix���3���1�㐥(�� ��9f��H��7���)�L:�_��pٓ��k����Ո�HDߪ�Q2��f�8��ǫ�3�7'4��X�,���4j�O���A�����r����N���P�/Q�7<_qM���Rn̾Nj��M�'��ŢwN�/ނ��03ngl��,yC��q����>H����f����*(���c��ʬ�e�*$��j����s�uj�U����CT�����)��YoMkࠨ�67H�r��Q�"�����2,-�����d�K\��BO���O�$�ϳx;�!零��m9�f_mxX������P����؄��x�B�||w��9����Խf�9j8���N�E���;�/eTA��e�yq��x�q5�S���Г��b҈��{W����w���3�ڂ�2t�R��8¹:R[����@/�'p��!o������Y6i[;E�k�~�joː��y����,?�v�W��L�P�#ϻ2�5r�~�!�st���Z}���W��FP�2�
I�ø�����쭩�i�^~��x!L"��\�f9����#�;�3<�1!�L�*-W@�;��#O*_�,\���u�R�Y-#��x�Ň���꼀���(3�#�)�&ΏR�&�PH֪ �t��'�ؚ׉=ϓ:*���{�y[\����Ԓ��M�����\H.1�����o����,�K[8����H�9-m:�h
�]�$���LrT�r&�Ùn.��D굚��C��$�4�@�m����t�Pޔ�y�z}dEasTb����Rn@M���?G��"�v4-%Ы�!��@���F<¾ �/���*E�3�)�5�;���>���	%����j����#�Ɇ�q�a�p9���� �#a�P�I���E;���H�8�g����U}!�j��"�U��e]%UJ�:ǯR�(lg���:Y�6H��9|\��D}6-"f
�{%&tP@++5٤ =,U+�O�5,}�@��y��j�����23JM�`��Fs7.s�������G}�R�w�B>^��:�%o����@��&�X ��#x�a���\Ԅ,4�em��õ`�L�����2,�M쒌R�!gir+*�X���o�u��<W�/"��&x6��]���A\�yG�+W
Z�4�`�:3d6�o�I�^ٙ5<�Z�gP�X���S�a2��@�_;U�Dܹ�����*e;�bq'�V�#l������@G[��f����)R�x�@�3�l0r��:p�����j1��^�v{��f��l#Qz�)��ӯ3}���|�4γo��]�z�d��Xp��hCto��Y�ۢ�pq�yZ+�XOս�)1�)�����"c	Χ�?���h*��C���]I��f���&��f��|�]�$��T^z�X�b�p�=�wRH�pϗ4���Y>��Ц�ŉd&�9Oz ��p�����ߪ_��Y^�vv����k���G�����&_�}�MK����'´���U�r�,������c���X*�C�H}�0f�t�Z竜g�6�5�N`�9S`�>�!�����9~�=�_` i�C�y' �L/�g�CR6�=�χ�Y�T~m�p��	��V�ګ}��F�y�.�Fǧ��i:����+���V������B	:�<5�=�r��j#RzDR�B,b�X�\��K��ݪ$"���пys��? 2�4ͫi�zwiW��ϩ��^t�uz��TNr���A��6���y8��eQ�8�_)SgTʭ%���^eܪ� N�\��t�=ܚu�'�C��t~x�9��v�5詢(�h�tq���wD�U�f�O�!�/�RCp��q"���K�-Qӭʜ����	�}t�G���;SnI�$�9�L��ƹҔ���'qN���._�2���M��A/*~�[�6?�TN�)�l.���_�-4��^3LF]:�o�!�R+џ�F�O[�S�T;\�DO������\��M�Qńhzʉ�x���3���/�m��^j
+�s�c���_4�*W�!!@
��~�s�GP�᷽֟{���?�;Z�WWr5
�����1A�t�(���!c���6$���`��L }b�E{Q3J�U���Ȍp�l�^�A��%���i�����HrPx3��:�/Ř�\Y�S�ߪ��b|�e��k���iA�8Rf�]���I->�e�d"F�'��O�xe|������X� ��*웺]�'��ͻ��a�d�H�����Gk�9^4	�u��� ��Я��H�_`1�O�0x�np�zIJTc�������j�~տ������G՗��"�E�G�La ��a���HJ�%������4��u��G��U��8�y~��N[.���r�`˾v�U� ��}.OuJu��b���o��CK�F��U�`�� �"A��G<����A_��H��۶ˤ�/��0mu�)#�5�N���'�:+���}���Ҵ1�4ʎj�_��w퉁�y�[H}p��Ȧ+P!���A?�ʓ��O�Rrzkom�;ѵ�S�\"����V(�7@-7ML�7=�Jc��B����ڻ���d2y?
���LP�=��=��G2)o��g�"T/j�"�L6��Pa%��� 
͞������㴾#�1zc�r׆ ���\�X��\�||bn)�.���ŋĄRT���*�>�Y�/y犝��'tU2��`�vr�9̚ux�*+��!�ՠ��ϫD*2�e���_��6�蕆�5<C��㜲���]�_��f��k ����͒O��K�*.w��y �����D�^�Xv��4�f�B�
D'^Viِ��NϔY�,��n�7��MM2a=��¢��#%��/�7�fw.u%!���+�>Pq-�'r�q��Ac�k��~f�����|'��!
�;�)����]�SW^u�T�_!��}o�����N�����ƭr���r�U�h���}S� +�[���s�X]�?���e�1	����wZ��v�*�σ���om�I�}��6��>r���S�ɏ7���)�ϓ��D]�I�p�a6� �#v�b.a��Pf�Y9�2	+�;(�y]?M�������KL[�ܶ�%�����<BTt���i�<�J y�]8;f�"���B}Taf,ܔ[���i���~YS��IL8$M��x�ܫۍ��驯�\^o���Qf�Ŏ�%]u���jy1�����E�=rx�x��'k�)L�m�d�Q+aF s��+Ӯ;eN��J8�n1�N�a]��u��K�m�uo��!��mշ�X��<­mE���\��%��2�>���LX(e`Ϟ�tj���\�,��8���kEt�q`�g"�2."�6�!L3_��E�m\	�}((�OC�,�z�6�C��#��*�e��\�G\�O�@l����gGz��7�eu�A���=����)۽t���/N�ȾA�p$���HVU<g�����4��Y��d2~
4��|�ctZ�D��?�����c\X��e.��~]T����4}�ɂq;��h6��^��B��w4%��e�2ur��H�/��+����d�ISǀND���hOM-���f��Sz�{!L߄詵�������I��
=��^#?R6Qo�6����J�N8����r~��>�	X��"�1���}���S
�%J E�I�CaT��)��(�o�X	$K�#�:3?<I�<��7��h��7�0�c��V��~�Fl֜w2�h�s"�����2��,>��w�'�k9�΍���4kv��P��9v4����a�tRB
s�
�B8�@��J�ыR�W8&�޴���q�ZG�%#����M�J�����s�ѣ�T"����B��r"Qp����!fj��ў��*?�>��RU,4�����="���Թ�/\�̪�X�m�͈��Ѷ��ZsJm�0#V�=q���E@W�)��m��E"�v�P�t2ha3!�����B-XN�۞�]\ #i2mw(*�h��'̃7'ca�U �U��Ц����� �.�k,|�ֈ�����m @�%Mw��w,����G-?6�q��;������PՀ㿡�O�5�ibݽ�blxL,�0���f�Y����Z�{�C�����@�	L��Y�������%�w�qѾv߹K sR�M-v#�N�)HQu�^�t%;rzڶJ~�HZBf>�jb��~?���C����0��hW��`�~ȃ!*);��]�L���pPq5�Lr������Y�V��J�I��~��lCW� q8뮽��C�7m���0���~��Ev)�h�9�P���P�j5�t��e�&�=؁b7�4�m���f��J^E�e-�jb�у�m��V�̺k�<��k!v%yi�7���C759�%�(�=���e����$��o��n�OZGvu�c��AΡ
���Ｅ�5��̙&i��<���O�Z�Q �D�$���cH���х�3.����g�l��+�bL÷�(�ÄUF҈�h�����xj��OU.�S��K���a{%9���u��_��ᷜ�I.?��؟���3�`�~owXF��R�MWd"�
���"}�����72JEӥ���m�y��Pi*H���LHq�.5%O�yP������a�EH�\�GP����t�@�����t޷>da�86�5����h�&�'����9�����"&}{.# �st0M����N.��a�$F؄����� �6)�}���MO� ��^����e��/�+��������V;���,I�'XV�[�I��A/j�U�D�*
��[�3�`��>�3�>+oI�r�FX9q� 1�:�o ��=�r&H�Б��L�(^���MDjy׽m2,�(х������O?���/�FLݎ�T �UXx������4��S@�B=�9Պ��B�N��]���z�g��W�e���͝�5!�$5�%8H�ܦ��5���t��	���e��'8o�f�E�uo\F��.��`mGa� �	r�u�5%5qQ��h�Z���,F�沄r#lQo��f���>=�a��&c7dӆ"��g�kń���Ҙ�d{E������'����&�0�;�Z5��h��Q�/*��{�H�n>�S���u����\6ǍݵR]�_�8B�>�s/f� q�:�����QN������t��󡪥r��1I.$��m��BU��/aU�Z���y������C��(�O��@�P�hD�#�`�#Jo�w=��ar�˫��8�a��踙��-oT��utN�̦|v)A��X\ (�Pp��l�%�,~M� L*�u(� �,�����q:k�Ky����&���7�?�*�8 ���m��}W�>t*�%r�/�r���X�����z���Kш1��Gu����k�ӷ��~�GPH��;E����w�cS	���o� u���E'�yCW�)���M��-<O���f�NT�z�ѓI�45ܬ3*��_�����i���F��L��,�b���G,2� ����|"�kSj$!���G��MSu,a�1�#��D��|t)�* ���|�G�0�mR��M�Y�{�S:jGZ�dTf�Ai�V܁�u@R��_	$e'#��q6��ݲ���W��_������8Z��1���1���n��#�X��%��~�T)sׇ!oxb��B�ϬY١������b��>�:����o>���� 0#`��F�<1hLz��풬�y��#�3H��K0D�'[)Ñ~2��.��:I�Y�J77�Fړ�0����>���O#�UjW?�����Q�W!�Jū��O\,u�2����)��ʬ�p~�K$���q����vʽQXޡt?���j��	���\�m?	L)�J�1����-�l������.������k�A\�iq�����ߍ�TFy�0�����i���(���+rU+h���}��B��P1Sخ�ه#jR������_�yq�T� T���s���M��:Dϗ1��Yt�d��C�Q��)R�z�vM���-�l=?�槤�IҒN��ų��8c��l���^>&$w�T�.I<ԚJ)h�nl0�Ux��ib���[�h���!I���]ks�0�n!­��vxsF�?sX��>\}�LuI\���J}��쇕f�Z@�Ղ��"����0���
R�(7}E,���.� �����>)���{��=`�2��쯳��ri�K��� ���p���/�TS�E��U̻��Z5B���Jœ}�N�ܩ?�Ŵ�t,߄������Lz�ڼ˧�B��?�Ϗ���#;Z�V��"� ��q��XΥ�~��BD*��Vq�R�5���F6�~Ce���֎xہM���ݥ^!���*,���yM�d|��A��8x����S6�Âg���&+[?M�X�PX�{�e$�=b>��p9e�u����{�=V_�KW���������`$�4ҍ^r����rVrȠ>�6������:��=֧ö6 �S}�_�-K��A�L�|�mX ��Z;r�t��[��2���?���ےZ�e�B]�k�ğ��C;MU���}�E\��;3���bP���߂��D+f�ٗe�q�[�wK��x ��YJ:��
�v�&�ͭQ�"�����Hț$'C^��"�xj��C�M����k��	��K��99��q0{9��{\����O<��b��L�j$�Cs�Z�~�ivC�*�#��9�g�D2���>�7�vn�%JD8��`��b9^,���R�� Z�D�_p���OȊ{�'sxFކ�0qifeA���p��*\�����~���
������Q��\Rn[&�]��a��.�^t�_hM >,Jw��o	��۬���+z��� �u�u4�NSL������&�NQE��p��Y:%cVeM�@mc�7[dz��E��>����$ד*ds����=Ahru��%��1K�?�=�Jo��|'{'����$ϕ�X����)(xv��V�t0�F�qaD��hOh��LGi���0uA!6�l��6�F:^)�ݰ�m�ZC��-D�s�a��hBF|*E^����������\;��֦j���mް�v��:戎��<e��N#�Lg�\��[�� �On�L L(G'�dɖSGO''v����g`0�� {k�F)�1�H��@��;N�$�r�����U��<R�]/<cm��N��,ț��e�j@�d�����	i+�<�aF-��c��
���:��;�'�;"��u=��J%8H�F�\������w'H�#j΅')�U���A��4���(�{^���E��'WeY�&�2�� ΰ�p">}��g�B�hz���R�{}/���g����pS[�ʺT\�R�n �9��t����*�זR<1��.���-��F�R���BG����C�j��ِ8�i(6��I�v�l�ԅdۘR���u�^:��Rvej4��q
kZ.(���9����w�&�T�%����γ}P8�D6v��X�<�=��F6�K�W��5%���y�������3�1��R���[��<5��k)"'�{���tJ>~�&��x� r�ASU��(1:����V]l� '<�`D�����
?�l�?�X�#�9�7���*��Bd:�n���ZaRXj���Z� 5=9!/j`s�I���{?ؼ�@�e��=�����yp̨S�XlZ7�L���(��f&N�'Ӽ�iRO3* ���ǽ��ʲAKA#Va�A��]Rb�	~X��m�(����ס/4���=��������,7��C�g���>w�f��=	ڑ�F����Pd��K�hKG�)����� �x����+Υڱ.�Az; ܛ�#�7��@�"/�!�.ky�S;�U��b}s��q$yU��[its�?�Dxe��z��k�4O��in�� ���<�>K,Q�quwAiFt��]Ӥ>��!?:���-ꦕ�YEw8o) N���܋y+�e���h'�I�y�]
rH?=�� ���>@ v�-�_4)��oq��i��z����x�	�=�:)[W�E��Ǫ ��O~���H���}�nHl2?�~��5Î7X�%��\�β���<�o��E��D�_�ٹ�hY�ƿϜ�IŮ��|R���_���B}e=�RF{�~_�(W�J�<�>�GaQ$
��H��T�3v��u��MG�T���V+Q�J��ޔǹ�[������*'�iET�!���9J8���.5<(c�К]C0G�#@�2@��'�|�>�C��W�� �=���u��؈�����('��v���v���n����+��c'T�Ϡ��نv*3g��O��;��yې&��� �n ʿx|s�z�(�z^OLr��k˃x������ޫ�Q�	��P3c�XN�f=��t�_b�m�Nؕ�UC���oq���j�H*jXJ'zp���f��G�CW��=�Զ|-W�����$Z!�?�v��O)�`گ���x�O�"��	�3|7��9�ة��G$� �[��oY�pP��}v����2��I��uFj��1L){�������v��ف�;�}'�EU�3��]�sh�I��e�p��DM�*��,��A�4yQ���W�EPZ�����͋���t �\�x���!!^g����>H-���駂��Μ��WbP�^�D�B����c���4)�9&6L��5�
�e�i�mzyԤ�$C~*��$��j6�U��n�����*�n��Ż,�K�HB�ѻ4��h< ��z��g[W>��.S��(��YP/�`�������V*)~����G�-l�U0�*�&�Jؓ��o��n{��2�LpQ�TKL�'��-���A��>�]��L��ڒ��]W��Rn>9�7c��Ҫ��F�'�i��,���̄�=��,�f���~C�G:-�ax�sg;0��]d�N�Ye�C覚-���~�%��-��U����T�D䙩(d\<�,[��3�����88�_	%���u(`T��r<p1d\J2�6Dv�7�.��'Awa�gQ[��oK/rᶓ�`��g�2.���Ux�i>@��l$GE����\ex�.��l�3�����~��M�7q�!ϣ��=;8���|,u��+�]�fiL(��J�&djm�B�s)X|� �P�����)�^2s���S�^�P@��[b�5vm�HkGɓ�d�*��gX%� ����|����=��w؁8�t�9���nX��m/Z�MQ�m�n�X!��U�#P=�n�D����v5�\��$Q�}��YU�5���n�?b�U�����]��Q��$IN�_��X��� țW��ͨ�x{� ]<�\j�U)�q(+��t� � ���cA�>?���I��,�X���8I:2�v���������i#�ۖ���S�2� E4w8GM���|������q]e�0�S�PsUIn�X���kv����
�����\�;�EY\���Ȥ������x�Qݜ��B��_�C���a2������8��v(5� 1��\yH��sX"��&vx��$oW
/��,.Qڕg�)ZW���n��0/��̍��_�E�R�~�
1�
�
w�>��!#Zq���HA2�7�������A԰��$/�(j�'ü�_�3y����v5b:������PȬӅT��c\�6�ՏGv��G%U'Q��=�5�S��̃�,���E��o+�B���3��8Ed%�!�Ks��_ͱӖE�Zn�H6����N{8ǅ�q�p.>Z���F���S��}l(م�ґ'�� ���<�I��L�޺�ޘ��\�ʐ��ɿ�b%mL\y�(kݘh7 dZW��N�*�H7�A.���#�_������Ļ^}ҩN�V7;�IDK��E�m���?���ַ=G�!�I&��B�-��E�-�l���5K$B�<�d�%�Ds�F]N��~	�ޒȕ
�d܅��Φ
B�d�Ab���<�ʣ6�"���)U 'vm�{�[ľ��HA":ԛG���'������5B�E%jN�EO�D��y��ٙ�Ig9��OJW%��:p�
ɟ�!��C*
j�M�i�ǰ�|��1z��'d���$mt�a��Ov������`y5�2�]H݁�����2|��M-S[��7����OW
�y#I����
�HQYr얩��e���fl��1f��r�\"�XԆ��t����e�������${�
ki>�j�V��f"���v,��t����""T?N�f.���O���.�(P�\B<>������H4z�I� �O�~�q�
_v���t��(��d%�S{�p��R	��u�ɦϏ��p�����V�\LdKH�!��Z�}̷i@+y�.6���Oob"�@��#�U����WJ��-3���`��8�a�2!fg�־�����c$���2��Q�Q����� U��V:�$�f@���H��~����x�(?G���ɰ�!�A���}H��Z�x��ѩ{��*=lS�ǧή��y��j3��(d긵�He:�,o����J2�|&���?���y��{jh"�m�P���ʡ�|T�`n��Z��2�F��"	�3�#Жk�.䱊cNQ���A���4�P�����J��j��`��IU�oo!��4~��Y;�>��14�L�C��4a��)�a���A^:�QQ�qd�a̸y�c�@����*Eʽ��Q�����Zs>
t��2��o�y��~ȭ�!%�_���c�.��<Γ�ӆ��򻝽���� V�Uw'��Ԡr{�d��V���4����
���0���)��㏖?�d�M`��4����Z:�I�����%T|&x,��0��*��ӛ�!��8-��5M�n9w?�D�)��d�U��~r�)$ٰ���<��@#o�\7�쫟/��6�)ڢ�Yvƥ#�WU�b�;FM�3�-��Wbc���z�.�6��a��̣�;�o��"_Г*t\���m�RG�{���;�����)��L���'
/���>i��(�����9�7Eͻ�}Pk��Wڈ��ttL�r��2c�vV'�fK�{Z�B��0�C*bv7Ю�0q�/�D ̴���f�_k�	y�Z⟁�͎�$u�3���N��K�(y3�@ S�N<0��:ުT�x���Ӝo�@*��a��a1j]��6�P�T�� ���|9��?��#��κ]�Q�J��+�oz���b�2������-[
.�41�$����]*-.�*\a�bP���lɢ�b�	��V�ٹ���^�}?>�Y��)!=V�!��*�V֊���S�ϙ��vF��|�z�~�e�3MD���,E�Ӑ����'��,�Ӆ���� ��5[ޞy}�ٚ/Q'���p>��W�/�/ ���Jm������uԍ�b�*$�Tq�����:)px����CEsz�W{(O��e�Tߥ�>�Z�l8O��0��I�Z��y�����?�8��K��������3*�,���%��B{�!�5���W�h��%Y�z������}�����Ԝ�Bg��Y�rC>�z����[h�&�ǡJj�W\t�^���a������q������%ݫ�xi���?���-�����Z���Q\�/T���z��i�t�\��%�F5wF��~N643�P�:���hp`	d�JH����o#�>��k�ȶ�zQxɸ��\�����;nl;��ITT���Z�7��A����lU�Ϩ=��v�1W�N���|�=�^�!�V�1�Ƙ�-~�p�!����p��F�3d@�������� ���Fv9e�"-��ny�I2������[����s�΄'��i��T���j�L��>ek��a �=\��X�G//���b�#���bj��|��h���W1��*5~�b�r�8�����Vz���1`r5�JH������>=�z�9��o�ij���^��|a����-�c�O?,0���O{���Α����|�G���T�9SF&��"��!��Y0�cY���qT�^ґ=��-(hi@@O���Mεo��u2��܂hj]�X��
�I�_&��� >r�k������ِ�tXi�vr2D�!���IU��.��N�{������t"ilw8��_�:�~�1�I�Ղ�{��ھ� m/��{Տ'e��-j�&I��S��%�٣`�2��,AM6�	�m;�o��"%� ����@�W�%���M�z1Y3L棭�pe�c�1G��6�h/T{�����������{�;��\�2��0��1<������l�!Ȥ.����N�;7o�Z���{{��J��n�,,�{��7
;E��2�;��GPp���s�/vȒd��W���K8�_�:��l��IYujrp"���2ރJ8���W�/���E��H��@��];�S�L��]��m�KP}�q��m��JY��s*��PtQ��
<~�y�bx��:;�K��O�ԔSl�s0d�ã*�w�a������z�2Ǣ�E69�J`y H?��Ɍ�֩3����^�Cc�/tfh5rZfz�3�)�]��!?*w�_�%��T�ӡ+v���)b��� �ì�I��s��a���ۑ`CO0;����7ǭ���kL�>cӴ)�Zv�h�"�����&��,��8�6�j�U�u�J���/V��p���|�"(QDz���S��mg�88�hTfn_ϔ�]�+��x�5�v+}z��Z��(��A�u�C[N�w?R>�Z�]Uh��܅,��7���y��>C�ׄP/��@�Ka�x�"bq��W�N�Le��ߥ��C����J��~��z*f�z2P`�{aа�ٰKNF{�ٌ�R��N�,A����g�vS�c**�F��W@��,��9��h �MSr
��. D/2��PL� �5Γ0
�V�Q`eʼ�����r�>����X�����;8n�O>���D�oE��iW�I2"T	�iWO8��G%]ސ���p
���� �3xz)�k��<B���DQ�Q�w�O߽���T#��L���j���J5qH�����Ĺ�Vw�K3�\��ը�R��[��-J}�w�����R�F��@f�v<(Jˢ�����X��YMO<h���d����Y�^l�ܯ��߰�����o��i
��(C��v~#��Lm�N���>�V��ڐ���e{���"z��@�zb�ȡY&3KQ����I����n�!.����I� �J�C^%'������Y�$c�bX̾�pN�s����S�=8w"����7\o�#�5�u�N�Sy򚎶�*�;@t�ձI��!��b_z��)S��Tj���{�V|%f�{��hW����0�d����f�G��tǒ� ��k�{nM��������b�¦������D��Q�1�n��/�u8�� �G^�5����;�O��ҙ��l���J-�e��FXFM'?d
D087Ȏ��x@���X<��7����Dg4���G�1��6c�Mi���T�폻K��fN�ؾ%�M��h̘;\�Y��)�9�}c�g�W�J�:���<䝸�M.�L��V�A�"&]��x��Z^NB�C(ī��_���YF�/��I��:�[~#Pݟ3�u�XC��VnOvX�@�x}��2���}M���v�Ti#�2%�U� ���8NB|m4���SCxM��A�?V~=��N]�	�1��9J��~��[�t�mi�Ԙc�ö�9�Ȑ�*|Ɓ-���^�����\���
��0���cK���W�8��ѝ�<�R�N��|�́i����:9&������?�LT|PNnj��fj�K�fX�L��a�+vbC#�cF�i�x��f�gP�8k\l�2���9Ύ1hѯ��;�<�a#���zV�:\!~�%=C��裦N8ֺ���0����6ne�V)��� ����Rz�HT+,Uƚ��k�{e�r`C?��̬A$l5�@�R{~����^\wN���mb��j�ᙖ���0;y.�٬������~ٱIB3��se&���� 0~jǨ�R6F����%�R�3��-S��05@yݏ�3����e�D}�k��!�� �MЬKߐ�E�,����ٝ�ߜ\��{�v0ӫ� ��~cZ�.�h��� D�ZK�bv�7@ͣ� ���<3���IU�v���o�z��>��~� �DZA ��@�p˝,&��ʲ�mz��Lڨ�72v�~Bo���ZͳV^�G�ûC^Q�QJ`v��P���"^���y�W�U쥋�� �-��e�ض�����Z�f���	�h�*ÂC���ڝ��[W�Ɓ%u<;3a�1�&~"]ʫ�r�5lq��k�3��I�ϻ���bbg.�����Vp�QU`WB���榉)�@�+�W�}p��}@B[ �(Ļ䈋1iF�!�����Qo6E[��OK˷r*�b`�M~,���C���{�nϗ�\�g�>mj�7����W�:�{[h�n��JH��Y��JL��ϵ\mJ!rpA����;��?�ɹ��p����@9����`���H����h����B"��`{���)N��v��^�"�@�_X$4������B��!Ǿ� ;hC�'�Ѕ��x��[@m�k����"�s��Jqb�z*v)w���ɪB�^��z7���*��&@�-:Ö�����j��P�)i\I9W��۰�n@	g=�wj�af�<p�gN�l�$�G�;�&F~�ˤ\�Vil`�n0� Vo1�Te'������L�3�*-��ܓ�r� �����b�W��i�l���Dw� T���D7V�Fu[��%�L#� �)Z��]Z�Yd~�*�Z�b4Uu�9�d��痁5Lk��]*-�D�)�η��t4�֫Wy�^@�P��J�(T%e�����#m�3�`�oq�w��K�{�K���D����9�U��Iׇl�5
^�n��+�H���*�"����I�˳w��1��]����s����h���i�jo�K|��k�%#�kdE� p��O��
Ê��-)�qriC�_�O18���7��Fqu[��)�W:�y��_#�EkG�h��v��[f���[ԙ+��F��&�|�X!��}��M��K��.\��Q��󵕊%���l���o ��x�jb�����q�p!O����u��*d�R^R�,g��[��������ͷ4%���1���Hi�<YTѯ;bf��������Kt��?� ��5��B_���¥����ӿ^���x���2�Y�tI�Y���O�c��C�,�[�!���c�y�g���o��x��hH}�\ =�@ʭS�jDU?�)��u�]��tT�t�ŇA_�R�gg��g
��~�8��� ����&�4G���[]��U�;tA����x�*�H��M`�B+�o���CR�C�pe�l�M����#���������n��=*�T��M�`~����H +P��<�mVca�ں�2�$�L5?��@�"�A01J��B7��ɚ�(4X��fҾ�j���_a`�wj/�	l:�?�X���ﭠ'��e{L�im웚K �R���W��@>�D1�'`d��eF&��X��YI!�q��zj�S5|�純�;%�~�<�)iD�wh�ݾ[j�K>��
F/o7;h�������4�{*�Z��^�A�7U`Yp��ܳ/��l�]�#�X�;R�y�.wڜ�{�p.�����|��8��!�g����h��r�tA�iE�#ȳ�������~[���� ��$��2g̾�,�
u��엮��v!��s����O'H��}��9n��I�2?佭-P`8��{�� �߿�|��fhoQ& m>P��.��f�&���P[׽�+�N���)��3�q�P�R͗�3�2`�R���N?I���?bL���|��w��.}xR�[��g�I�d�/�-�t�Ʒ�C�^��}1�7$�g��
�`��(������_c#Q��:?�z	!�ob�&Q��&����{x�; !qۀ^N�q�e ��2���{�p���[�$cr�
%�ZK+�3S��l�.�wP��8���\��]�AEEu��y���Y$]~Mmļ��ڋ>i8�|J|Q�;ђ'�Jgȥ���i����q=�O�M�%̂%T����$x��*��mN��W(�Tzd\�Tz��cA�/���Y�ȸa�ҒuKQ#�T��sB���=��|�Bm>I�t��|��|��wr)+�"L	.�=�U�в2�$u��\���'��}���ņǯ;Ȳs�wk?tV�WI)1�)��Бn��e�M\����Is+�k�3�9��OV&�1-yc�
W��E��wD����f ��"������P�PJ^i)��r�[KY :�����%��N(�#`Ѕ��0M�64�
����-�LrX�a���+�΋ޯR��I&@	�Q ��C�o.9O��vC�k-}��O����v4ѓ��e l�)���R���'��i��k�VT�d�o���G���J��CGy�Uz�ɳ�M55(��%�S�Xx2��p��5q�hU3ڕ�^�}�~�s@�frM��]$E�Q��F ȡ`}3�'��ׂ�Y��':�e��cd��[�ذn��4Ѹ��P�䫒�n�=��Pb������t�^٨p'��3��0C����(r�IM�sV_X�`�9D�t\�����aD藋�2̛� 3�B�/&���2�D��;:�~f`��.5y��%�ٴ�I<s�x��t��i�Yl������u����8o�t�gFΣ�e�C���&q��[��"������X9��[��)Hs�?�,Y;6�G�T}�&��i����v��wP�~�Zn�pl�N�;�ْ\�m���=ۏ�Yrꁤ!��C\����Rt����cy�h��S��R��R����d0-���VG$
�@�=�h��0�ڞ��j��楆<=J��y��Hb[���qq.\�����l�.� � fL���S��Jk�]j�a�99l~
>��E`p�lMG2�~��!Nj���Z�ܮv�+s@�:�͡C}a÷�yt��[��3���ђ��y�^��
V��H��>s�n@q)Ǉ�s�XU�[�_�d�^�}HD����p�2U�Gb��א,�$ڈp�LC����rI��R=�ӄ׃��ym�-��~τ��`a�gq]�n��v�7 6w���+>~P��=��\��q|��"�ɒ�I�r-pz�ʰ�nN�������V�7�|��S����*��&9��;v� ��WB3[�ʿ�����b�x�|~�>��䆀$��<2x٥�J��CղAU����.�}M,�"ԫ� Bf
��h���ڃh�p
h���"x�x;r$͔���	����e�!�\�OK?��>iQDs����p�"���2H��[��E�&�J�a�_묥�O�z�4_���Vҭ�X����d�.>�PpS�s��{q��<j �92��+܍rm�,7/���'���� ���剞�;+.z%6c��F�n�?$��-i��':.��ᡱ#⏁X���!T�`��[b���ZD������F���J�y���.��Jd�EAGZ�d���<+,`�-��BUQ˨(�@X'�4t㊫�e�h� fj�=ĸ��~R^ݮ�V�]R�5e/U@����1��Y_�I7A���LS0"5,�Q�e�V�� z8��]��#�rڏ�o��u_Q� -�����!��{���)�*���,xA����t2��A��	b�/�G��6Q��?yJe���I|rח� $E�cU[r������n;�4��$���5�qi`|�K��>������Wc �x�w/c�{��O�R�*��#'��CYƘHƅ�7߰>��"�����B��7����ގ�ۜ�H�wH�ԯ���sƥ����Q��`߷�%���3TQ�-�\��7��`#�?7��z�!x�-�>�Fr��Q蛹��x��˼��@r�5S�Y���P�ux�.����ٜ���#�-%�lr���$�^^�V��~�E�k�}w��U&�����-}i����5F��.�F��!'e��A��N�p�����Ro���Y��ϫ�
m�?����T�Y
?�9�T���>�:$Eh=���>c��O��SQ�"�pN�o�N��N{'#=�����&z��8^]�מ"�n���A���H�Q ��FD����	έ8��ݣ����y<x)1�o�~���,�	T�m�^S��v�M��?.���-��E�<N���o��d1ІZ�P-lr�k���b��T�g��|R��.V�7�_D؄s(�G	G��o 4�Qd�I ��Ү㗂�(u�N�HnK�_��	+3-b_�I.�*a�n6�� �7�['�E��'���{����?�#o�/P;�x�;W�,�C2��T=��0cYM/���J��.��z^5��C7�7ae�d��XǤ�"���} 'ϻ�5 �궺|�w�DL� �W8c�e��
��[�� �x�����+�В�Hӗ��>*���C�	j=xJ�H�G�Ӎ��cs�=����	����vƈ����9\�_���+�w����igD��7�Y�݅��̺���H���QNJ�}�x��Y���p��002�"�`���*���4}�@�B���2����͘�8�d��C�{ڨ�F2�#���1ڿ(/r��ܼ[J�~i�~.���/�a~c\!����"�����ˏ�9��c�"�P�fHY6	�B�,�wւ_u��)wN2�~��Df�=n�m���ߩ�Ft�l"��5��8��ȫ%�xj�趆6p����h��?f.J�&1i�̬�����'.�`�fK��V � �C�	5r�I�� U$xE�>��f(}f_�,Dbx�a����Z.j&�
Th
�⁛�/�F�!~UWM!�:��s%�`(�\e�|�	�װ�?Q��_0�k.�+lxD�M9��r�|���q���S��5F��x�~;{c�UP{����N�6�/g�L��4�}+F+#�OPQ�L䏢z�f� ��I����`��Ϻ\�����D�o���ږ��8���۳J�$�na�������(?ԋH��>@b�	���8��PU&*(m�[n�*�����h����[���$�@�v���ž��Ӭ�.��l,7��H��j��L�U�h��Y��qO�3�|�Ep�B�,&�t�öG�<���W^S�&6V��{��F�1pIf��40R�y�W\���LNJ;@<NΚ���F��-�"����~M-�X��Or�a�#`�9z��*mZ�<�n�9�'�u�B���R�"��R��i3G�T k@V!����[(MuoKˡU�W��:���a�:���p2�VmW��O����Sw��A�/wgoBKZ�'�7ĵ5Vw�(ObegA��9^���I0�*I�`��6�d������ުՊ��H2�xR��~hf�ה�>v�r�>����6�Q��3�������d�R��p�;�v ���FvL�I�I�� `�W��f���)Ќ�jgsu��1���
N��rv��K� ����*���#���Yz�����c�E.#])�%ͨ��{)�ʹ@&T-XrZ�Ji�&���^�<��n�������\�
{��zƜ�/���_~�Vr�M�Cѡ����e{��>m:�����4+�mgzVI��o�m;B���z�\N�=o���2�gJ�ֹH�|.�k;���E,��e{���_�]��;m�V!�4ɛ�� �X�ӯ��3m@�6X�AYBr��s�L�l�'� X�Lʟ�����Ƕ����3{�n�t)U��?GСت�:T�X��E+���>8>;��i$�m�r����^�o*�7�`�=��������;�c�f�<�����Liy�`MHi���a w��l�Do���=G/A��-n���I3����DǣG����B�/]lv1��ɯ�7����<9�
`���\Wk=���5 ���*�SR�nE�fAŒY=����V�]/��&��W!��g��San��X'��Y<���Y�nX�k6D@������"&
���(\��h�mz�g�Vr����g�z�^��%^�_��������o!�,=z�^��cs5�^��ʅ�\0%�)+����l�~4��-^�t-�s�/�B�@���o��OgP�p���m�;���x�BRi���m��!��0v�F1�t:�M�r�+��
H�o��j�9/��]W�.����\�+�R}���H��<����a\m���L/���,d\�V|�1\2�9�>ڧ���}g��t�����^7'j�%�����θ�̺�Q��?�|+�Y[}j�b8?�ٟ�ZQ�N[vw:#dKn����Z�� �|TJ:���G���6����9Yb'�9�Vڠ2�?��-��C�� �����QC����i���%��m�U@t`D��.��\Z,�K9�k~g�e\po�ARC'��_?�y��D`(��)�a b��3���XУ��9E��.(��h��QW�@P�x;�����I:{$�2�ڮj��3���'���C��oQ�0Q�]��4�1���0i+:b^źT9I���7�$	�T�O�)҂��OP$sU\Y�u��"���z����^��\z�E8R��;ϳ�A�>]7uI���@�H�5A{����rG6����9��d�I�A�I>�� b6:(cOH�k�P��a㮂��� D=�M��9�)���q��_�#J��Z�ϑ��B"�c;�.�sx���w�VB��`G�4��Н�)�
�vW�U{G\�ի�-[�,N�%C�����[��$�~�� D/�bp02�u?!z1�({底S>�����C��tCJ��Occ�i`���#��x��Gh�xT6g�{D_��?�֧�D�����n���0�����[S?���b&��*q0���"x��)��7�5�U�A'��0>���V��y ��V��Ӫ6s��H���Y�aX&E� >Ra�A�s��=z��Е�V���ӛ4�0�D�N��Q�$BC}��o��lL�0�f�����~pGB��v2��)p���z吏��+�L������@��#k��6p��1��֝-E�`)8J���B�CEK�8�?���|<��J$A�;�V�PXJ�0����u՞Y!4u�YP+3��>������5�̃�`s�EPm�t�]���1��uuJѬ�CE2���ٛ\~�*z��;d�mt=�R�ę�O�gMm�eK���H4V�D:��*�$�3�Z��و0J�4�P�ǋ�:�#&��H�$c��M[���^�za��{��PG�?>�z��Cx%O�&�14r�#!Z�'L�k#>�g�`������j9@�+tY��Z�O")j'�l*]�Ӳ�� y��W�&n�ct��W#��R"LCy^&�[48YB������Y+��ͳR_O>�x]m�Z��y�9x�&D1H�^��L�:Q�߭�n{����^�$$�:JD�;م�.~�Wbf%��>k���[�n�4m���L����:3Xc?I2FQ�&�R 9��������� �OZv�wں���*�Ō"�BL���ǎ>�����͟�d�Hb�R�[`|�k7t���%���R�=�7�����'L�ͯ��"�z���&!� ���eA\,�"�Ew��<��E����9���	ۖ��T+���LM��0K؈���OT�Y76�-�Qtč�e&���{�=�d-�d��mHtc}=\o)�� O�����u�0�^�]���21K��葌��4�`�n��^��4��VW�̕�e����JQ)��BzWr��+"�mch�B#�9�P+1������?h�N�PãEH�:a�Oٙ�*�O~8��t�Vi�ۂ�RH�`ҵ2��s�shR�ݡ�c9��rz}�|m������ߐ�C�&���*�I/��З{�Z?_�V|���������# WT�U��++E��v1!\>c�n����p�l�x�k6����I��~��{Q7�n�~�]�����V�s��%S<�HɐI;�����Dw��� �ΰ�w<���(�dd�AftG����6�#���=�ycw�'��*QQ@[�%�y���B���_�JO(�]��|A*�j�����ژ���(���[���,0��8��$B�M�<1H#~O$�97Ӹ&����e��*�����P�'r�'���o�!c[�/�,��]��E�V�x�,��]��Ї���k㥆r߭e�s�ST��ᕲ�\��N��v�
}GZ�w.�G���������g4�I��/`X���������8�\��$F�̚���g[
���K����r<3�WQ\g�c $V���?�NȀ�^���J=��X�y�&Z�(�	hp�	?���!�;���\,��7�~ISNe.;[�ld����<�wF��U��v#��-�T�5K�����AwI0� �;��n����u=��
��� Rݬ�23e���9z2���O֧��r:�)<�)��I�$��hJ�c����t*)��R�\"͠���6��S�s��������Qu���;s���������taz8ї"A�&(8�!�В�z�sZn����B��nV!���������çz�[�C���F.�R���H�W��G{����R�r貟�����/)t�΁�Ę���_]f�!���ѿ�%"uh��|R��b;���EE���t�]j�ܠ��F,?�	ڢ���[�Q��HZ��R��|�k��FD�s��K��k�ӵ]�%�2��������K�x��ڍ�W6��bA�����{���׮���Q(n��a�W)7ҾN7�x��Pg�����DS]_S$D@Ҽz������+�\qɼ��(�>�-^�#8qtl�༱E�Uv�Wg|�{�B����� �A�*����@���ݚ�f�V�2�t`&آK�D�Ʀ�PhX��1� ?`�B��#Ԝ�5�JK��xJ-�CL�Qq8��A36�hc� 8ɫ�p���O�
��EyqT!�cL���te1�:�!D��2� ��?pz�K��Hs��rd�t�E�hbzq��K�r�ņ�_��ۺ��P��n�_��B�Q����a�5éRFm�+�b��^Ƴ�8f`�`�p�,�l��DL����U�`Q�_��[����Qq�2�u��яF��3�ћs�{۱vJ�"K.�h�"
�!�Fl����Gk�Vh���Q
v�+_.��u��x>,N��9���6Y�!��%� ��C�yQٵ3��7[�%1x}��L-�� t�
Dɓ��u62	7!�M3��������i�giwQ�VĚ��m�����G;��>�iZ�F�Q{��hI�u��PЂ']H]���.z#~�!�gn�B�K!���L�Z�����)o�Í�%��[���W���^�s$䦷*0M��잣F���	e���o����"��ׅ5C�e��T_}{����(�P�.�?�[���Y�'���~��?6�XE�7�]:��S�us�<'l�(R�x8�XĽ�c�Jq���ʏ�J/wؙ\�M���
	!��؜:���A�
�y%���"��U6�j,�3a%!?��wb��E1<u�jC0_o��ڈ2���ٺ��@*ۄ��*��#��B�tP�Z�����sj�s���A�f����aB�]dO�k��]��i+9`s5�V��3Ŧb��e��Y�_�sw�@̬HӬ�\3R:������'�/��$U4� �����	�
rG�	�g�̰G�ZS~ �zO���:t�3n��Y�m�������"l��i&�1A鎳Pl�q3�:�E�y<��*��ct�`_�]%lo9 ����@ʢ˷ɀ0�~Q�n�S5Q���3YF��_z��j�Q���z�IDǚ����dK0�d2��q�Ix�g�ŕ�`t��d$]"���6������#?6�%'�I���_�`�d1�H��O�b����#_|��C��n^x��gI���Z9�~)���q"�� ��i0x��J�� h�B��BoL��6j~���̥~0Q�x֍V�v-,kcq��1��7���(H��`#�@�ڊ����Wq�ps~0����ږ��0��"0ޭky�ؼM㲾����yq���
,=v���͝����9�h�Aˌ��H����PY���3���FqM��I#����'2��۲Uy/��D��O�������U�n߽��dG���*�kWl�L6G'YW�'�^0�[sŠĸxbWduڃ�-���e��x��� ��KqmR(���\Уor=t� 
Bi~���Qc{�@�5 �kI��)5.>�vg)-R�k�LX���ˁ)j��?�ݶ�?;�J{�ɝ�c���Y�g����͢�\-M���=5%��bM\k��7�����]EǓf���>&�#0��˹l ��T�j��J��h�dU�;�� z�ԫZ�%�)>.���\GC�"� 5�!��q�v��Z/��n��MǄ!|�.�N�a�x�o�y�B��>�>s�z�Ѱ,sqx�f�z�<���fA��9�O�>p%���|G����n�T�Ox��7m�z[�jX�|�+�=G_)0�����&D"��3'������Y��0��.��)|4D�%8u�2`n�)�/��'�o.?�z����ڰZ��:�UMu,t�K�"Y\��#x����Tb��vq�Η��!�מR�TM3'8`���76�R��e%n�_s]Z`A6ք�U`���|����^W���!L�x3s�'���g��`j�l�۔�[�S{�DW�ad���cc�5������#`$��y6�f[$��Ki>��F��W\\Bդ�Ӝ"�Iy��������+Y���VqDZ2G�u`�k[�yI���[v=N�����w�H���#�j���]�}�����'d5��Eؤ�$7���d���2����}�����n���d����)���N�3�"�������]�-�9���_�oẊϽw�MU3�v-]�r������u\���X� ��B�=ڦT|7
�[�b:J����Q�\}�mI�nM��1i�J�}���u$E%��5�Ԃ��pCз:�}��a�oK�'�y�]ׂ�����$�8�"On8��=
y5��m�JO$B�P�rSؐ�ٓY��k#μu L�i~�;���\7ߠ�8J}/X+Y�O����I8�����[J�g_1Z1��"4�Q�x낛�K9��4������K�G���������Z��k��׀��Lx�!��3n'�!7�	g䄥��m���b���K���t�O���9K �P�Ů!��;�����G�� �ώr�@0���=��^戒���?Wο��|��Gk5Nf�͠�W���:@D }"�D�-�ƀ~ԓ���-^xlZ��[�WM�h�"�ޱ=r�ИA�%Uwj.C
��1�	c�A,�W�C��=�;t���ܚY� q� �Nؒ�Yv@�W�eQ�f�bb�9�mB� ���
u��de9N@��_��;�����l�������w��*;��7��$���-q�7�ȉ�ږ)Mf1�OT��s�W1�U�R=U�����|�MW##�1�����k~��6�eU���ϜJ��}D����b3ۄq��TI��;B��ص�<�/�~a3"/��M�tIw��,�S|eY�+.T�V�p�rY��'�c@�
�a����&vE�ɉ}A#:?���o�y� ���u)�C��4��*�]�\	�c#}���[s}W4�}���GE��n<��є0�Mn�+O��b�h���w�ԍ^uU������'�6�6�T8^�p����r����.`���s�]���"�ޥO�{���s��H�Xt]k���:L�f��3����q�(��-ٺ�=6�&�R���p lhb �"ǂ�Λ�*։��GD�S"�Q�o�ee�"���v���f�؞B��16r�d$�;m7��ó��$iۭ#��(b�$��(����햸a�`P��?xd���>8�3K��E
�!�>挦��eן��w�MP�r��,rq��X� �U��o|`������*_'�����Z�4�)ǣ{Q�vga��I�=K�k��?,�c@]�9��SW�q��1q���:x��z��.�:���R88�'Xx3�גV׼8C��ֿ���U�����
'�|7�It�:�J��@�k�l�p ��/���Ć�-F�4g�rI��U�o���Jj��W���cS%�Ct`��s[�tȼ��h ��Z�	���+_�i�i��+h�� r�T�a��/t��&೛%������l��M"���!��J%��Do��H9N�k�.t�-RȃW=��rqr~� �Q�<�V��w����.޿.xy����>/��o�xE'ܽ�VὋѓc�����ż�f�!R(mŴ�Q-~�"��T�����H�D�<������9>�Zf��K�%^w�8�>�����o{��a�ǝ��5����K�,�52>�� V	��$�l��Oh恏����B��+E��xu��4%�E��D�^JA�ڹ,�Ȳ�?Pr��������\����}m�6��O!1i�~L &��sPx�/�j=��g�:��"����^E�\�[.����[��9�!21�('岼)�>%6���
Slה�:���fK��/����u��A[S|	�6#Q��X��	�f����+�rf��>KTNEL�z�G�˼��U$���&��FxY}�8��*�Y6��?��|w��S���qh:mikǠ�NHЕ3[��~�Q7�^���ъ���JzmU��k0����1=)u�uy���*`>���5�j0��Ul�*;]����ř�Q�t~_'��)��nH�R�2�W"�?bxs�K�������+YV�F�����ǬS"*�"�{����;�}�M�Ԣ�)� �f/YJ�y��&�몿CdZ���V�l����U� �>����R
��6�+B��(<ݳ�p���ZNgw��]g�q��:���U2~NH�6C���h�-�eR�����F���$ď<�V��g��#�;���m\�� �R$���D���ىpx�+H��WE��u�����..?�;��fmvd�{p��`��Kc��}���C[��aU�u&�SGu�%�?Oa���� ��w�T�GB�^3g��Ӷ5���O����@:V��*�y�2��ZoǵҀJ�A��K0��|�	J"���&
O�Q�ɲ0�@�w����N/�36y:-a��~`	���"~��|�л���S|r���z̧ �(�\cL�8Fpa���&�D�Th0���~X��h-��IY�xb�	�O�L�V�>�D�z�����?E��9�"��P��r�4����f2��Ѳ�RD֫wC�4gZ�H��s���qY8��Qg`�7���|
>[��;�Q������T�Sey�{v:��$ע��׎.�ʿ%o�"�0�B`�Z��&qH�m�*2T� #G��i>������1�9���˲FD��[�h{wtHkpwgKVZ��� u�5�SƬ񅺻��I�Q�a��*�h���Rѹs�wnWw�^�A���U@�5�$�7�r�D1EF�3]l�qp�ª���N���mbʞ ����i(��;D
f,5�j�.ӳk��>�]s�0xָbzh�'q\U��_�Hc:^n����w�|��߿n2F��&#Qe������<m��Ӝ���D�C���1������L�֚�Rg���|к]�q�Q�d��� <5�X��U��eIȞa8���D�EA��;�wRM���u%W��E��ҹW��5�ȅs~	�V���D@���"\]���ع�X�� {���@��5���x- �U}�7����:�Զ��+�xY���D�NY�t�)H���U��piM���$)-����u���$?o,�l��ẵ��nk�Dɛ�g���ؗjفה���G1����0�K&��!~*�Z@��=Ȫ���O��Ft����	��l�^m|GHIj��[7r��H�	��	��r��w� �P�MU2��Ku����28.�V�e��1������l+��G�d��AJ�)Q��ͱVr����
�
wέ'U�����.s�oU����]s�3����?����;�s#�X�aSng�0n����i@=8�����J���?
��i�u�,���v5����s�*�%.�?T��cp9@��*?��>�Em%l�eG+"�������)��l�cJ���ى���@kߧӻb�>����I��s���<̒�Y�J���l]Z�͘j`4�]c߷l���tN�`R�*���v.�A��6zHh˝$�H�����+�.���5پ�Ά���$[��KZ��KJ`�\v���yD8n�����&����>c�PsOv�"�lR/Eԛ��*�U�;�+��D��2	U��}WD�v����T��ֲ�0��(��c��cu�#O��%lR��#��������@v��+���"��TR>��m�uz�/IJ�haV�9oj�|������Ϡ�|�q~�m��l��\o�k���E�^�Nމ�&T�'���7��7�_6�˥��"�$顬o��a�0r1�7�u(���~#���+ݝP9��؊+0�[���'Bz-�Ɏ9��VH�Bb�<���͂��] ��'z�/�%8ن���������PN�l/�=��� �"!�l��~f��r�|?�&��>>�z�W��[B��C�����j��#f�FRo��>��t0���t-��v~�^U�Ь�x��0�E���7$�%��Uj�%�=SGQ�h��u����'����c���+q��P�Z��0�僯|�a�ӣ��Je��mN�=�"�5�m ��^�˨��mۓ��&��st�n8�7O�͒�������2���s�
HO� qf����= �=3[<��{נ"^�����+��/�I�wU��98��A�\�O��ijt���b����Z"��hd�u�8E]��q�������j�������J+JL��2D��l�%&U�|�\�o�.��e�X?d��O}�D���j�DE�	x�M)(�9"��q�[/L%Bg���G�Zb��9%�5�O���z*��xaw��@��ma��ON�nHi�C����#F~��'��+�� �_�_y!�oC�-&h��f�k%��*=ʾ�M�����f i��/QL���'D[��>��O��s���Nƙ5QN;Ы@j� ��af+�p�rG�RI����E�,�O��DO�^��t�:��M��~=t�I���qv(�3N�[Y�z�8:OSiD�P�ٜ!��
�L�Y:�;O�F�綤�B�U(�^i��C���v�h��F?��se�uN�F�]Gܟ�>�����K�El�V����1M#1Njn,*,�n����A��7컽$�+��%�2�ì�9m����&�4�
�R6�T�G��м��� 3r���me`��x�`oׅ&T�=�÷�pŉ	�T�[ޠjU`��	��>�os�0�6��^�9%"X}��m�|�[��KLY\qT��ӹG�*�k ٓ��&;�Qؕ���%r�yf�����'�^B�|�O$Ň;��$_�9#�o*���6!��@ޢ=;3�Q�I.�&^���}f�Za������u���v_�7a}��"��O��r��<;o�&�@�n�u�Vxu[���4A����P�ԙ^c�C;�I�r��:��Q�F�������� :�v�5���u��)��	�O�SO��ҭ�R�I	L��s���|��N���� y�Ͻ�`�9&����tv���'#&_�7�ЕIՆ��J����R/��C�.Ԡ��.�n�`dU���T)0���b�x�[�������`��	��<�����;3α��o��o��ΏFm[N�9�d)W'���z�J}Ã]	Z���-�Hgu�ˡ"�-\�=�����=/C�O*�w�{�RU�� �1��ӻ6��G*����bqhN@Q<;��y���ȭq��ḓ-���x�c6t��Ē=����v��8�l��Y�t;U9�t�^贻!�5�D�X�elD��g0N�H �VPt�Y�D�(��(��٧x�z7�+�Bj7�\y�c\Ӻ3J�LO3J%�~H@?My)�3�n�4�cDZ9מd�s5'��P�5f���Ϫ/�"?�aa �O!�*�1�p�^s��s&��YK�:C�=U�+��L�M�1�eA)�خA���`U��ޏ��I�ZK��qx�H��J>�ֶ�|�d�xFWvwP��
.2�|' c��~`S�M���V�	�^z�{Ld�[�1�Hj�z E�K],�Q}��٢�d�;T��ϢR�⠿óʇ�ܛ�HH���\D���3�c��U��T/?��3���ǫHѿ:�Q#��yL݆.Q ��7付*�՘�#O�>li ����
� �
6�I0��)'�{���2���3J�0	A��`k���OK�&6��iX6Y#�B�zː#
Q=���3v��͔�5stA�"������O>j�#{�L)��)�A7{w�BԞ|�F���	z����q�������ډ�SeAc1.ךZ7jB��-�m �"W�@[�4X\�o�^"��@-��8����YA�������p:g�y�=��_}���5x��������2ã��$ܟ�	��F��Q� @T�]�����C�h|��@�v�$ݭ/�
��pg�<ral ��;o`!�ݡ��{H�Фqr�i:Տ��F3���I�����\y�[��zɒ���1=��G#}�(?T���љr�+�Cz��`�C(8�o|��`�t��ny��@���#9<(qdnB=y٧1�xhx#*�>�w�5���ؕg;A�KMzI���;U�S�<.��IF�r�G�q��68��L��v�>��;�� 7#�xϩEyNC��3�.��\��&j�YX{�mH�O+m��)�������4v>��:ؘD�-�|�S��k��3+�����57���V�/q��ѭGB�ӌ���%�o��%%_���r���>�r����'�v����
ύ]H��7�����RUս����~L�*�����B��e��:��������D֛����od��%z�x�-�B���WΡ]L[!Jx`N�}���?��8�dF@wY�@I�� �B�S���1�=�9�s)�ደ���a���YN��mCYQ�p_�Eo��ʤI�� �ߐ&�U��O^�pe��|���+t�d�m�*��*��e��Ko��E�)�^�59>�^�3t�/�_��8���gl��礛rᬃ5Σ�1i��[��UX�4Tᝆ�:�F� �@�҅|j�Q�G��T����|�e�.�]I_�,t ���j�]^�*Hy.�z�Q�v�V �͋��Y�P�w��>�lb�^|���Fd�ˤF�,na�Tr�?S��i�����!��4?���,��q̄���&T#�<4
Ksj��:
xi�pѴOpCw��5�0�������VI��5�[����+�Tl�����TJ;C#"��a����D��0iI2�@�9�$�#�aPa]5f�f_���v՘�+F�k~DV���l]|ls�Y�=���j=�r��f�Sc6�<Ty;��/�nE�L1M�����{wgl���(�\��;�=$ˋ����b�ËUb�P/4i7<g���9cxOET�c@읯0��Ώ����۵n�cu�A�}��j�3F,g�UPR�h'�N�,�����/�4�l�wS�ϸ����K5����)D�ը`0`d_��I��hUk�b��!;	x�K0;&���&�6H���U�������Z"�fj肒�A˖��`_[���+}�����o��#� +�؝�������;�v��C�L������m���97	@ꯍ��q���5/�� ���#���a��Ż�+I荹��yc�%�a3�z�ХLޥ��j��>�ӰA�z���9vͼ��I� �eym7�S#_:J�,��FY+H�x�}�&���s2:�nL��דd���cj���HZ�x��* !�C$�Y(�FJZi��@��2�㛜~��i��G�p��B��E��^���Lw(6z�ͩ�������a ��:)c�cߕ�F}3�`{ƴSZ��,%�i�	Fm��S�7�
z�]P9��R�~�P9z�E\J�_����4X�T{�X�`��a�����bMi����٤�f/X��IEʲޔ��)���������rf����z�d�P�h4<_�F��	e�b�Y?�gj	���7��x�I�Z�s��Ga��O(M�e�Q���r���4�^�u������7�d� [@kK-��*JT�_շ7�8��,�X��83ǚ{&ڱ�9������l�D��i%Ӗ����k�0[�0L`�Zr���\��Xp�k#s��+���S���͵|�-�W8L��V����
�k��"��a�7�k���5/�ʢ���&�䅯d<�
�4r�R�0��7�HPj�m-ZDE������+��A�qC�3��\,)��m�4Qb�:�ؑ��T���]��&����ۚ=#ɼ:�2��aޯu�Z�Y��=3q[��� jRcB���+����nI`<���f��Mxl��,�:XQ��Xpp�a�����ʐO\U�#�1X�Q��J�0TC�X1��?�24�;�zT�+v�P��ԉ��Xqt �o��+1�q�}�d���E�p�(��t
��m1=����t��#X�6P*��.he�-��h�)�4��@��)�T"��6"VB�sN(��m���q{@!07�1Y�dm?��Wч�﷔Y��Vr�����b�^CH,?�#��,ş\ⳂB+�$Ӊ�b#o6��b#�\S��YW��OW������91�
<���`���Y�K�v�ubEp���x��Z���xL�cHO�Ox?V��8��]���KN ��s�*cȠ�7>t��k��Ag�����5��k�����}yܣ�1d��Q[�T�!/�gWHM�\g�=(�������`�6&��o�oΊH���[���$y�*� |Ak]�jnFU�"�x^���cޫ:h�,8�$� 0K��Nxu�Ffْ�D���w� �n�qE6!��fqX��W�r�,YJ�cq��b��ڱEG��]Np1$�c��-�%C�����e�(a�a�߇m��_}�hŌ:G��4vM�V$S;��%�T9}�󱄼]�ƿ��[d�/A�݄Y�4�@�a,��@�]��1��J8��P�nw|q���?�/��F�4���D�
�&"���4;W���� o-�6�h��!��`�"^M�,� R�V#f8|����4}���(O�Pa������O,�*M����bੈ���F�V6)�ެju���X�ٶ '�
���Ah��<+�� ��r��Y��cY���,[^�J�GQ�`݇E����͹X7P���7#�B�"�_�33u������dZI(��03�����8��Y�܂K"�L��3��DG'%�2�
-g�ZF�-�I(Ο��ڡR4���U��aԎ��3{�%Ώ+�XT�ײ�X٘C=��)�a��@'���y��̦[6����P%�&9�����n]�;-�(���%�3a&&���m��	F�"U��fES����r�	�*4ɖ�J *�F'��Nd!���bg-4�"������'�'z����Y�&��"�-E�ax�����'��J$�/g�߉�h ����wv����_��� ��D���Q<X��ܖ1m�-�����!���}_IK:�L��d1�:�����I��};��8��n{ ���B�KƤ_ %�V\�N�/�&o{�q��$�#i�tnf��]�����׊��]{n��{=�^����)8�$=���~'p9X@���o����Y�1E�aΦ�~���O��w������Y����.e*d���Ʃ�Z�Y�&آ��6wy
�~4����kپ����Ak��l:?.��g�h@ь*��>J1���0�6�E%�ߟ .Am)�')|HH�#��5 QJ���[f�LUI�߆�����o�v2Ϟp��U�_�M�������A���¬zKr�0��Z#�$��1c������r�j	�K|W_�`<�+�a+v�xx",�QY�x#���qK��)D��,Hj�ܯ �F�*j*N֎�n�h�!�)�z���y�(��,�)�(+�2؍gOA�e�:!St�0s[��K�nQ�-MՍO��ϲI��3ӑ*�D����>�V����pK��4K�Dl�kǎd�8Ȼ�Y����>Q�6��
N��T��0Jɛ��|{ ;Z�`/��:r�U��-���{[ԩ��)0��(F9���9�,��Cu`���"�D��1� �����nK�
�n��J}�g9)D�w���ȷ����g�"��^�j���U;�~8��4�	R����6� e�뎔b��8?��m��FB9�F_�d6�^���B�F6�ͳ�Îb/[U'��d[�q�6Ǔ}7�cq�������/���D���j����wI��Lmԋ�q�!y�T��h`��k�Yn��-�����H��������1��@e�E����ΫGpN������D�fz����X_�y.��D�;h�=⺦�j[,PΓ�A�f����n�E�^�I盟��ݡ���m�h;`�%�<,5	
��jǿ�7G����#)&z=]C�cpvY/�Y/��/�ڬc޽�a*=g�Y:%���Ug�*m��~��@W�}Q�4�5v�AD�C�*�D>�\�~�N��9�L���C���
2�^�5�P��2�`f�:�> �����7"d~��x��@A���NGFy����JR]��9:<\�g�CH��47R��d�2h9���J`� �nbd�-��ќ�;�.��$9�<S�%���b��O3@�P�I�>�4�q��	}6�� ���NP�K�D�Id|{��&�+?�IG�c�AW0/�P�=O w��S���qJ5�J����xP*�j�!4���Q���&&��s�BY@#�x�oW�r�v=[�+���@3�5
Q�
�&�$�Oǝ�p��l��8�&C�O�����\�Y�e��װ�w�!<I�܌������3?�j?;� 6R��-h��L��u ,��<��r���%��z��\�.����."��$C��H�Ӊ�`�2�v�f��р�\Y�YD���)�5ʡS������US�P���*:��8�T�~7���F*r�W�Ö2�%�"&�L��#�bd< 7U�⭹J���@a,�ʭ�D��-8��_���:�c.N�HW�;�q,&��=�â���:�,�G�g)��������e���X�L����?�H#bB��8����򰰼�gDS
��*�R�1p�Z��������\r�ixd�*�c�L��?ߐ�>FV%��Xb'�z�;u�fyvؤ�e�?*//V볏�!�ȕ_j�����,��s��� �1P�eYh�R�Ks��;��!�
o�_9�H�a���n�⡡R6%���m���&a;���ք2l�y�]I��e ��̖]��5{�{\��e��y�(BjC��z�3�AKL+�����VPj/��ҍ��Ѿ#�hĐ>[�H�Z�R���8��r#��:x^�l�4���������(�0	����?h?y	��s�t�V��;�����ڹd�]���˥/�X��Y���Z���+�uf�'�e'����RA��ܹ�{���%��a"�T��Xw����#���ͷ�"VIDrg�.=R£lk�.��t�6�3C��|	r9�4����� ]b���u��Vw��ϔ�ЗɆ����J��!4l�XF℩�Q�[ҹ�'8ƭ����5G"��_\�����>G�-��~�����r�M��pqKa�tC��_��`W�U�]e.S�u��)��ߝ[n�+��Q��h�b�/7�ȕf�h�{��ZGB��_yh�S� hɼpu'ZL�e9
���X�:�fԗ�!��O�Vq7��0�h�4��b�;�ˇ/m|��ES2��D`��?҅�ğC?Qv�d������-���'�V@��a;��@n >��d�j����<5���4��fQ[��6d��/Rs��j P���-R|:l�)o0�W�A���-:��Z��T�����w��J�R�騄��&����-%2(B0J�����8i�K��Z�id�s2�s���N<�M3����MCG�B����,V�(N��2�</�6I�dM��&� R7#�Z_�2?U(	����VQz���/�ݻ��&��y�4E= ��_�$��ߣ1��&�+5�t��bE�gL*!ʖ�����ޡ���y���5`˭CUpԝa�a.<�R!�h �;�I'8"��{�FP�R���U.�D^�Ǒ�xR��NmH_�G��_�dN�Տmk���w؜��|Z�J�@��%�*��Ǣ���>����U��;~��|�1�Pn��eT�=R��a���&��Z�+��p�" �����jϙ����[�~�S� a��22fx����YJA��d<f��Ѿ�qS22rڲr`�uji�\��q
���!઺/������<{�e�P\" s�L���w��s�J�a��/�ts�7����K4"�>��������6������)��;����m���zJ��I����U����(sa�b�:��&A�*A��y+�������� `3��jg-��	�ov� ]Lȸ�f����NO�~(�,o]�$7�������|�c��l�Չϣ͒�!=�m�1�nOE��#�tD��\�d!�bU��]o�1G@�Y�
���o|��ޅtz���a����tT$��~d���b��S�h2$��U���'���:5�2=�Sm�������N�inUk�`UG��"h_TH���J��OiL!R*j�V���h�����?��㘄߇��B�X��V�j�w�h��R�9,�,:��A�D��b ̲�mD+.^3^��,I]���Q���z1#�:������~���skP���uBS���}7b~�,ݲ`b����9@g���`͟ ����� Vɦ�3�Y�"̣�n���[�hS�4�{,���A���l�I��^M�F�s�P��'���=2l?�<	� ��D%�������q?���;Q��S�E}X�u�'t�R���e	��x43��IpPݵuR�\33{|��S �3��5j��z҉�SDI�8���3��25�W,B�y����̿�/o��k��K����l��i�y4G��F���-��IqGnĻFh��Z�C3���.�����y����GXh]#T�t��Ne}�'�̑!�@|<���!	-���m�������~��O��-��o��1O�i{$kp|�p���H��g��|u���A$H*���ۨ��7�7.*��ļ"",�&����i��o�'�jZ���}��{~���E�+&E���1	�8X�G05O �qb�)�O'hN侶FuCf�65.�phk�*��c`;�҆���pg�W�����dt���W�z��lE�y����3�Q8��U"�#G���,maaw��^94��D�yN������B�wh_Ax�83�F�a���I `R�`��6���3��鏨�C��ivnlx9��Qߓ��vO�;��G���i]� 3��ꀅ @7`'�k�?��DU��@;O��,|�����6n�MoC�j�ǮW��I.�{g	�KmF�Lㄢ�����P���
�Fa�ʊ��X�v����q�Co�o����6���H��5���U����4����Ks��X�
i�(б�i16�r�N�A�0l��������l�C��eg;lvQ�8�'��z�Zz&_�H��-�t`bb)�x�ΕAm7a���<��,	x:.�N<U*{���xT����n����;/��H�������2�l*��h����\�5b���D`z��.�S�d|[
U���S��U�.�]�5D��x�-Kz/+1�kL�Mj��4�j?�,�����������K���F$��Չ�_b�N�A�,"%V=��u�Jd4��r�`Sǵ=�v�SǢGՀ�`6���2��s���8_SgQ�H�ڈ����"�埨F��T�?X�kvT��~���O��� �����(�u]D�GL�bǱ�ȶP��ա���*�yMvar�8����ӱ-up���&#�-�LS����('K�v�c�������R~�a��D�Y�A��u��z��/"�Ї��'�������ٻ��6�T�j8�,g�4O���'��{���4s�?h��G�@�o)���Y"
�c�s�����m��r:=��G��!�Ik��4w���P���ȳ�'���?�/h�K��դZd��X�v�m#�@��WY]�q4�a�Ed�#�t��m"B�V���]/S�g�j���7��k��g��2c5%ݲuv2f�cv(�G�;P���ք* c�z�TR�5�	���f~$6	):��qL�$�k%�Ɔ_�1ʫ���q�y��l�b��2A2)�� (F�����+z���ǜ��Yټ/y1������և>~4[�1� ��ݟ�6�X���6�1e��L7����jY���ا~T��y���~d�3}�H�t �sx�ײ$�����} �cCH ��jx9u�r���)]����u�t[%l��ِ��3��|r��/l�]:&ٮm�F�[�1NUKQ�%�oi�7
h��D�?%�cx���&k�7i���6�S���<��5��K��xy�����6-ò��K�W��>�bl�9��~� �q���� P�hb����T��`}�mT�T
N^AХ�ܗ�Fb^N�� oخ�z2�s����6��h[*^���隳�+N�j�+�ek�x�|a>@�ձ�p�� ބw�{Hͯ�I�ՓvOB���6�
k�U7ߛ��C�U��T�o7Yu��,�|�0�X�xт���)�	n���������^X�_煲YL&ձ!�p�'�T-%᜘��h�����~�N���̀r}�,�Y#��l!��Y^�M�y)
��m�R/�v��� u<��r៿��/]rr�^��=�nWpy����	f:�&�(��j.?qu\��XVh7�!�	X�:��f�b0���o�7�I,�_N������wf�|"m�yB!9��!�i������Jkم�R;ue��i�\�|�>������f�BbG�ʱ�{p�A��q8=|��a�Cy� �룹r���
N�j���@�y�����t/�����&0]ׅ�m͓�v����UM`��
+k�O�#h(t�����B�X?8q�%�F�ʞC���jW����{��O�1�L�?%�`��=w�����4�������R\�PXW���@CE��(���K�pk�O褋���vh^��߭���7¿��FwY,s�e�<��I�Ԑu&�<:c�҉n�D��	�-�V瘛��xf��nW,���3�V�[�X&�x/c*;k����0(��y}M$��cg�[�E�|�y�� �������gb�oQ���>�iC��AwS������#���~tW �t�*�Q��R@�'`�¯6f�)o���-�'��B�*����24�+f��b�?ۄ�*�-����2I^����_�V�� �M�[����5���j�t�Hr�LN���$�?m�E�A����#�J�I1ɺ�D�k:�j%�'�W��W&�%���{O�h����������G��{o����j��0�CYL��g�r������ V��}��t�n~*�P���vL�g��!�r�vQ)5^9F�'�1]���	ҿ��ء���&0��2S�� 
���'F�.wC|�ς����J7�/]��8_���;�`��4����*�Zj ��)����l�h��$�ʔ�4V!�;ჰ���ZN�����r7+D�W�v�[�^8����Ux�8� �˞^�D�fL������6k�\i���q�	������h�D+�G��+��L��Y�L�A_w��Rx�'�v�W-ǀH�`��� *�46�&2g)�t"1h��!�����Ҝ�"��@����"�n��I�hWS� ����w4��n�IרH�.6����^��9l��2�w7�0:z7��/�M�h2��/d�^�����N̾�U�6%�"��y6�pݕ0��y��Ws1���&M�[���ܘF�p�i�p;�iV~x������`�%��b5�)�I�>4)Մv�gl��+����ظ:�vTCԚQ��U��+��\�y�5Dj6S=c|#4��(���q�o�w
��]�ҩ5l���R��d��4Nُ]�_�����SU�\K�M$~������'��s���P��Uũ�N83��6F��J?"�X7e�\��G�B�U/uJ���p��c]�4�;��̈��~	���k��ǎ�f2H��� b>�o.��[��a��?B?��0�=Gn�2�m0%=K����|p��E��@e~�G�p�*z����T��f�Y�*��O0��+_LI]��Wɝ��K�_n�6��
�S�iΏi�
�(�#����CTk��okr�k7�Q����b"�B�L��*��t.p�[�h�p���L|PQ��̗`교�˻$2��n�LP)�� ��Ch<?���y����u�a�.-=ܽ��+��bN�s���?b�
lJj�a�P�Ck[v�|K��|��A����VJC9����i8>}�n<��:3��+ǻ�C��A�'�z�/|��K��|M��Yc���Ԥ YA��zk#��f�%���PF;琖����fz�%FQ�s��ra�8� N��@?�B(����k�)�y�M��sv��Y����G;���e�@�dH�/B�����Nߵ��K�����=��Z�*=��3]t�X�n�n�Hg�����0��-�.����"N����Q_1�!��*i�A*�1V��i�_h�^B�Xr���p=�x*�U�s���:ZB�0��&�Vp'8����/tI|W�߷�-oj2a~%?�[�[šR�Y>��e\ϏeZ ��!Rz�P|��k��V��Ý�fJ־#-q;�ߩ�*����3{��Ľ����p�y�f���c3�y�J��V��|l��V��*h���ƻr��w�@><��.��V�W/b��Jj66[T�l��L��ye)�ԠT29�����]B�XW���t�z�f��y��k�%b�8z��~~G+	le� �$W�ί��9�Y,��g��M��1A��2
����
�z��*0�e��gwk��Y9��|��w��icU'-h�M�u0�3�a��3#9�G�i�}��>g�>K��97i8���`��(�_�y�(3�x��\>�񛮹򯋇��P��� -�����W��,,i����6\P���o?c�!�RUM���\� .�`��_V���@YIY�$��'��-��V�_�]Ti��<���ޣ�ַ��)�����ܼ�K��q&2'������?�E�8�t���X.�ܕp}5�L�x1{ }8��@�
eP�f����8�E��)��M�����R�7��Run�lQ��_�Xâ�诿+V�luk��.Ɍ�E����Q
�wj��y��n��T"ݨ>� ;��L69z�Xۇ#+WO����Zf+5�1�{���P₫���r��t�D���q�_~^��*��	�~~�&��3�	$�C$4%x���귈g0�r��	h"+����ޑC9g$ącF����'J1ϙ}�����`R�b�w�N��"h�VC�&�A�G��B� �&�ހ���1�]��7D(lP��������d�>���?�Ր�~Ti�j����p�O��&�Io�D���O}�x��y��VF�x��M/�`~�ؓ��Z!u�ǩ���*�������sr'F%:%�LI�Ɇ���/K���j�4[
ʺ����+���P���C2�*�X�����Kw�Ō��q�˂��T���mb�ւ��~�~ߝb.�Ӄ奐�I��?���-��+�m���Җ*o���9 (L%f�8���qԹPwQ�$�:|-*��y�'�c�m@�zD����Iܾ46
�F��/V�+6>T��G';ğHXN_�ؓwÛLը�Z�w�#���xt!�6&$��4��Ù@�F��N��L6_�G�ZG��b�%d���I����$��-x"�#yJ��EX�H����O�V����J����.A8c;�R���N�qbW���/�1�K4U_�M0�2"8��S�/\�����F ��QP,��4I|�|v-�-���)\z�5�i�fsv��SOS����4� X���tu�BNy�є�=�>��C���
/_-�4�O�
4��*��Y�US���i�ң=!��Kh��Kvt��m�hw�ц��PS$�$��s�}wM�Ga3�M����'+�s��aƥF����I�{ҭ,�Y��a������_��g5�Z���lZ��U�j��x �
��u3�-�ȯ�-}���t��P��jjਆi�r~���0�L��UR~]/��*��4:�,��4f"�ڏ)H���{VjRL��O�=�6�[�ų1Х��J�]%�ۊG� ��F������&=��[Nd�\�s����������(�b�*�}�g��Ҿ;�b�<C�a�l���	�һ�8^l�N���0LH�5i;:+�h;hYXBWw�*��Mq�	y=����{(W�?�����J�̓�Q!q�s�g�y��N� \O.�m%��Ve@���U��p��@�X������<r�[.�����J��v-�u�J��B�!�%DB��o���|��A�iT��KT:�ZH�~����������է/�+v�D?��k+Օ<��{��Ep���~���xUS�:2#�v��=4g�6Z���N�OԌ�t����C�����Ξ(� f��9��E��C��q�[ߐ��u&��̟>��Nxm�. �kX�ۈ�_<����;�%`�yB☄m<	U��͜�
ZF�*���GC3
���g�����$�Oi,�#���?.Ȯ��߶�U�z�|�Y�>�^A�՜���G��3��(�[��?��h��گ���p�yC@>6���?|�̟�i0U� ,�9k��c���=�kv�@V�� �"D�n�һ�c���grK�%��x��l ~�1�,�MB�k"�К)��-r"���'���d�rAt?wlj)�6v�w�к�2t�v���L����t��.����ir�F�o��P��s!CoxN�|>�Q����\�pA9N�i�7�ݶ#�$`z`�uf 3<ڣ<	�(��*QM��	? �,N���;�8( Y���v�[�cbφ��<#/-^�n�W�R�|���R��pd����bt��
Co3�I==�~K���Q:W��o��S�ADCx�����+����XX^)�.�����܁��� X<��j������� c��-Z�*]_��/�<�a/Q�� �Dԋ�н�Z�W
Jm��u�!����2m��O�MP�^�'��}�k[������MNp4�[՞��2ucm�0X�:�Jc#��p�����Y�XR,�d_c�ؙȵ�9 �M� �x1W=ꢇ�����������qIĎ�P���t`�˞6�����.�TC�N��&����+j 76������<�ԕs1��hrG�P��/�B�l�X	sAT�fK��N�c�4*��W�y�4l@�ge�Ő�ix��M�K:�72"���q%��H�����6�[N���β9�5i)ẀIR3���2]�VY&,���Q6�a��6����G�Ǣ
�4���b��0���cՉ�j�]J��.j?������D���-�,I9Q<�P�Z�&����I�w�bJDn���׵�R���a��>z+���+1"�B���^���o���}@(%4{-�g;��`|Ｅգ�L��uD�,S
Q��\�6u/ɏ�_5��gN�`�3�*��Y�5I��Yt�y���������/�N!�"��*�㛒]�0�A'�@�<��)��t8�<��X�j�@���t!��~�6����W���UL�*��C�}Z�����������������B�#c��@�`N'�\ҿXP�(_IAj�ZWu&�}Cv.> �Xn~�+�B*\����BV�vm���a���D+KߌLW%5��\�88�����f�"�s�?�Q�'�QXY�A@[��p���r��Bp��]a�S2�?�9�p#;L��������y_r���_�a��"ap��k�A��W��Ģ�s�["@�v�ߔT����b�t�I��6f�t�а�?y��A����+s����Tp�ۼ�h��`�K�C#�:�ė�|B��tV�Cj�N���s���@O���"C6T1|R�xwa"���^��EX�rP�h�4�/��s��hCk��J�!��� \���_�j�'���#��M͊N���ie�*e�<�ic�6�����\�u��
qxQ͝��y����C�(��
R/vX�F��ƹ�u�4���v��I�0�1�G�f�\�E�9��{���dH�)�f�|M?�j�:�-��TSR��y�Mn�%K�&v�}�;�1df�X�"i�MM�q'���1�9�H��
ޭ�R��W�:Q�ճ�r���-�y��� ��?��Ȁ[�г9��.��-�g�@4L�C�.�:K^��BEGOҵ��h��u8�-�\�������Fq:h������3��&��e��.������6�E��A�Ë��KDч���u%y�ɮ(q����f�6U�Ak)%PuK-7�|=5�v�@Y�����Ř�5�Vl��mu:��;75>���܂ԓh"�$ K�s���溠����<!�<Ok����jtȾ����������ĺ"���L.����V�N`<���J���|<A����_93��.�;\�ا�0ҩe�v2���:���:辖1	Ƚ'ԣw��"�G4�U��퐼D3�w�-�W<S�Z��3d��A�Cw�|�)��}�l�x1�R�:��9��G!Cȩ�V�e�j.eR�%b,�\��A�O)
}��0���g�NB��U��X�����r��(�P�� D Q�#�@����|XvD9No��S�g����.����DM�w��n�=b��:w��l�4y$�7�w�X�2�a�a�#!�mU�c�Z�n����Ӎ��	gT�%ô9Mް�8Y7k,�2CP?� C�a.�����?�*y䘀7⸱����Hr�n�n��eE�1&r���E̔�V3˳���,O�,�|e���v����x�
nY���^��7Ͽ���X�Dk]�v1���pG*��[z�R����y�@�a�u��|�U�dH�	��vS$.��P����3� x���v�ɔ�͈l'nLا���­\
r�Ҡ��?s��#L]^8����L����{��.6��R��B��9�Ŭ��NХlN�ζ���B������ZY�Q���%P֊���b��L@w�k��K�	!���#�	�x4C9T���_�Ϊ
�� �qݏ�S2W�飓��o-qF�b%���vU<mg����
q�m�N�!�W4�\lG�|�f�/E}$��u�mׯ*�(�xɈU�B�qN��rש������H�"�3ꢎ�ϩ��-3�< ˧���%D��#��#����(N����c�kAvվ(�C+&<�ߟ
ʅ��2���N�O$v�����\S���
Z=�U������.k���-�=������:(���mČ3�WȤϚ	<�ϼ������%{ؤɩص�eI�~~Z��7.����,5�Y,!��4R&K��	��5�]�uR-ت��O�z��pl/���ߡ�6)��ui
��ğ�`��wf�93���`m�t:�@((���u�0��;�DE�N��p-�|�u�mXOr�s�$��H땋��.I�b��Ө��O��� [@JH4��!�J���I��^S��5xL� ���~�zCZ�k��h�%i[����kj���������Id�A��X�Kt6|bs�`yBJ�LAj�ʹ��9�d���=�a��=�nͼ(�S�v�%�f�^l�rs�L>3HS�rw�r��rK�Ќj �>sqSә������Z�������h����%��O���h�F%��8���&c�W{,/�\�f�+{L�q*<�OE��T�c�"9ި �����=���u�뇱i�R��J�+}�cݠ��4<��m�7F#R/f��������B�����`Z�B�A̿��gV%T�6s��Rɷ�Y�B$��n2���h<;[��:�#ͪ�\'s3�����^3�	��*��B�v�b�:'�5�UAp/��r���6x�P�|���N��GP�(!��cb�g���db|%���f
����f����1�[U�:fԿ9x׉z+�)�@�&-�1vD��뚝{!��y0�1��o�����;�Oz���	O���~��N�H����a�d����!����*�z�S�GT�]�Jsb�
�]S�)�2u��#Ru깶IF_d�`,�N��b4�&aG�C�tI6P,��iX��X�m�L+��u����[I֢T}kPY��B�ȕ-W������#��p��"�����g�ʲ����%n�܉���%�G������
y�볱�YE"�F -���)���6����e�ו�\
}�ڏrR�0Q��ƅz����`��|�d�K��c���$����F��175l�/�����7��e,(�Z�a�0꽉؃S���&�C,�L�߁a�n������@�W ��[��U�Vm��g��}�t}6�����7Z��#����a6�!���� �x�����h��8��{U��֮}q�Ö�Og���d!y[`����*%�q �/��:HH���Q��x>�΍��:�#m1�b$�M�oD\�!�H��G �����]��JɣF�<E���S�Hb�{�V��
�?P���F���ɨ�IIAEwӼ',�����$!�v���Ԇ�V;U���\H �O��6u���vJ(�A���G� =ˠ}c>wG�H��zF�~���� �����Y��jW�z8ƞ��3ry��X��v�g�~�<q�Uw��[ve.���`j�E<�p��K��ISR;n�DL�Ié��2�Rf���¢�ٹ�x�u�e;���TQ�;|�1O�����3��W���A��+i�E�5��ܜc����_��PY� SP���j������9��N���+��-՘��6������9O#4����ˠͽa����Q�V
-�1��0z�ʑ.��@	�������e>��.Ŗ�����p�G�=�=�I릲����QJ=�R`�KO��	���0r���.ƻ�"���|���Ch�����R����p^�/
ɼGeL�Y=j���y<�X�,pS8�(�Al'�`?�Ȇ��r~|΁�{�z�G�D��R��0u`���h[��yJ)��.�Y�����x��
5�u���ɛfL��^O�Y�rTf�Ǚ�p6��b�T�1�	~�Zo�*�#���-��5xl!��ר�}�&~����Z�JM��h����:Px�V����D}�Tti���d�׈��W\�gV牗%7a�%��7@� ~>M�����$6���y3G��}&�3J�}k�\v5�<#�d�z��HI!;+�����P?�mM�ٔ_���+!��ec�䊯��z���R3R	[���FD��ߞ��Դ�Jgc��0~�����D>U�4�c�Fv��L�,<1M�ك� \*1�vd�3f�����!��^���ieܧ"����\[�.UD�[���$v�t~`����^1��˼iO� U}�X����5�}��7I�ɒ�Bj��Y�'2��P�����5%8q�4(.2��2@G�\��g�������&���Wn�Z�V��Db6+,�KU��f��ѤO�I?]����d=БY<�)�5�&�Q�4����zh��i�m��{���B]QD���z,5mR�|�XR ��F<�����k"�O �omi�̛BPE�w�PN-!�ut�-������aXW��Q��[�ZjITR"S�S�K!U�O�b�+Y�y�Z������r�?�jb*���((ctzm##�A�̧�?8N�Oa��@�D��O���&F�1޴5��KpIn��xf�h%?*���b]]�/�K�lQU|v�z��]lī�����Ye��x��푿�c\_fM]|�ҧ�f��'�f�s�{�!.HPt�It��tI��!��,���[���2�ˢ�O��D��U�ǆ�s%~�ϭ����.�S!s~�憷����u����Iȗ*�Y߶v!Q\�6���a�{�Vu�����7���"!8���D.������2!V�X��y������l��10a���)�<�4f�r��G�v5��D��.u(��+qU]���o��5���KO\.�FaTޟ(J5k�&��o����zL�3��Z)ămlH��|?��پU&�����N+� ?9�d_�A�������o�[�M�p��VH�S��oP7۵���_�|?�eO͙��qÔ^ru.�0FN�rO�T'��?<�R�wGK�{,F���פԟ�U�H'm=��ы�r��`�4ZC���W�9m��U7�Q�"X�
��s����z@k.0fn'����9t&�kueH)Ҋ`%��791�0��)w�Ӽh�CL��غ�R�]>n�Q���(���b��*�*��Bۄ��c�҇���/��)#��T�Xl�G��6�B�����V���L�����Bz��{f~���u#/$�*񞄈a^4�l�B�i�����,�fQ�U46��\�{���$5�� r�0��6�koU�0J�[�>���"�HC�aU\I3���d4�(7�4��"~� ��V=�@�&R@��Vp`�6ɥEM�	�Q�p="���%>�P�+�ܼ�l��P���4��;�㋟O<����ū�0P�-��0Di�Tu�F��v�g���'�5��%��ʦ��5�o���=���;6촙�`z�=�H���0�DÄ�^h�>uH�p�ʓ��Dw`���V3S)fg"���@ޗئ�E��"S��W�M�t��`��*o��W�N��-0O��w�Q�;l��U�x���ue���n��β�C<ޙ!�`���?1I����ސ����hſ_�t6�N�_�d�*a3rvA# ����f/��vW��Q�uC7��b �#�~�r�����ʤ�ؘ�ձPt�X�؏6T�5��i�tuq�h�z�2t�Dt몐�$҄4h��y��.XqmV$��
�DG\�A𾨟7!�KTЍ��+baPL��&���)�]��w�(�ی�O�LC�g���L�h`�9}@�9 �r>��� Zч��}/|���1�f%j���}DH��v?�+ߒM��6g�*ð%���.饿G:S�D��<���jAc�K���f2
z�C.W�_L6�`��em^[�7L4A"�:�b�*�%�����̙u�}^��	��}纼�~��l�X:~R{���,�M� ^�[�⸀k��oy��,Կm�X����P}�f�F�T��}��`�O4(�S�w�Br^��k����誔D���g�&��
�x�΃�lKȱZ���ڠRŴ��<�$�_HOSX�Yd�P3��~<'��]Msgꅺ����eo�y���{n�I�m�L�v:�V8GgW�1�ZۡY��	c�lwQ$,�X�t��keؾ���oG;��%���x�iCK�{D���";��:d�7���2��E��<,�z�K>
c�p`��XIata$j��s�xx �"~�n�}Wrيgd��UkǪ�.҆����p ��=�B(��:y�p�&W��t�t��1oKua�i8��d�L�m^P0�~��
����ۧ����yҚ����������*�@����~���������0
S�o=�dp��n��V.d�.��&���3�3��3��oI6�̊z�q�9/�Wϑ��<�y���c�U���51�f����7�l���)ms��ش���@���MP��7(��E��^��Z�#���Dgr��bB�k.����r��M�1�4���ߘ�`4)�q�G��e>\'`�М: 9���{�E�~0��`��ru³�9��j�����Ji��LoX�����bi��<mG��N�w�{Q�V�@���ͷn=��Y�<��Xz^Z��b��½��nL��O6�~�ٱ�50ƥg�"�V5i�����!4�&�N��YCS
�|]'Emq��B-�]��mp@d�ǂ���ϴ��f���2k��H.��A@�r�N/�S➟W�evEd[@&�-��(35�gaG4VE�t�[a���;��?W9��g�ѝ�7���m�_�f5�.���߶gȞ2.ZiXr.I���)J"�+��@M8��Y����P�5/�2��Ggk��\,���|�SlX/?n�3j� /���9m00�g�B����RSu�0$�$��?�V�d��!>���SZmg/���<t` �lm�<��X����Kɞ�̷����nM��1N�h6;������J�����z6hS��� ���Sc=n5=~B Ag��$���4��`a/=DW�)"3��Q�X����m�lߣn��*_y��%04@[��@6#�s����Y�j0�eu��v1�l}hry�r�a)D�p^DHU}qL�?3\o(�ݡBSqMc��V��|0aH��'�(&Ӄ��c�Fwk'�MB���S��g@A�f9S|r�yӓE�գ����T}$��̑Nd!��1"���@<nÊ9o�m�90�R�V��X���Ip�)<kI�%.��*3-�O�%����*����y	�˓^�^��o�w2F��y�}g�_�l}.�e����u��k#`���$lP�1R:��6-�{��s��?%١S9�r��o�uHg��p:E
+�u��/hI֠�+D�2~�D�IƘӿ�.k�r�����Z��5�F�#���]x:R|��-޹�Ds��4��ө�hQj��,R� ��f��z�DxΌ�% ;����ҭ9�$	��-�>
n��ХZ*�,Ӧ�����d�bR.�%:�~C�x4*��R �c�mP���JK�y�E;c�;1~ST�ʉ� �$a��P�ցP^G�^^��ܹ~��l��G)�It��J�b`Ͼ�ƜM#��Īg�-�ϧ��R̯��w�3p��;
�re�|�͔D��Z���َҹя��^�(��/0���닷��]�Xn��f�"�D�m%M\��R���7~6���0�4�TB1�S��'��J�|y���p �n�Rq��is�|do��:��]2�/��u3u���eh�����ZP۔u�M�G6Q烝��&��`�/H���E����! �E5%�U�kpf-X����K��Fֵ����T���!�\�h;��#�F��~���4���6V)��������w{�6E]Xg&��Nj�m|��S؂Q�ںޖ��+0�Ͼ�"�/�.5j�TmEe��v��&E���G��_��0W��]h�+J��%yY(Y������Pիed�Vr�Z�R7�lNb�<�f���v�X����Q���/,��q����UIn�0�����f�DVg�_��?I:/z��r�r&@^6.6�tt�@����L�}WE�]����z�Rc�#6���
!CL�o��d.���\,yhlN�����q�1R��vru���HG���X_����f�"�;��,х;o�D�1���8+��Xr_�ӓ�搙r.Cl%WQTgV�]aZ*K'�!k�@'�����i�0+7��ҡ�Nʷz��:�m�}?$�/3(�H?���뗧3�ͧ�}��Ֆ��ǫ��Ͽ �t3�B**���o9�v_〩p~5� ���l��cs��ǆ��x@�bގ���[�YJl$jy&��{iV��!��\�5D�J!���"�H��za��f�D���P��@�`���)�2kw֑���b�.N� ��\Ky�����N°$�*�B��k����QN8��'���n��ͨ�͞ψoj]��3��X�z=_��ꩋ/֨�O�Ԅ���`��wW�Ԧ��M�Y�(Y�9�I���A�_�ʂ��&��e��7�6���Bݭ��Y& ��\��{]�SKB��I��_h�ZI�`���kmƵ9Z���p=I5�p} R[5d)!�!sE1"�jѷÐ�&��s<��8r��j �hH>�*�)��&������T",���@����?�&����z#ٝ�2�TZ���L�5!�k�C&JԻ��|�`�Q���pQ����J\R[T�0P�-�:ra]�i�Exr�9�P'�V�jk��QF\�ݝ����gͨR��ț�m?Sх�)�t�s�I�CR��*V����R�%�>�����Ⳇc:k��$Y����:����ӕ;PÏ�LF��|d_�H�}E��+ú��C
;M#=#�񱈄@�2�V�]�>�0{��U��ʾ	���3�d��*�*�T3|�x�T1*V��z#�\��aSmXd�E�X��6D�o�Q�Λ+/N�h�LY��X<}�k����JI8��N�����L�+(������,2��߱Q�-z���	a�M"0�j^�<��sL\x�G5�?JFh�w�˜i��+j>h�Y^!��p���
M^�;ܼ����]�A��[�I�?�}��K�8@�֑��(�.KzL���Ȥ�t��X-Ok����QI7_8l?�|�uj�H�R��ԇ)V�ⶇP$2r�q��ꢶ��c�i��~�����-F����>:O\���y�%���A%/�� wD��p*޴���	�^�n�H�t'���clW>��p�3��}+�����i07�31Xf9���Y�xͥ�b�v1������3�vZI�/�C�^t�)�<�E|ay�ZX�쐣��W�� uc������k� �rnqs�Jg�ʨ��G�n�܀2 �~}����&�=;E��֋�7TѦѡwD��F�_���a���8�q��X�����&{��4>�T+�3�zg�&4��fh{�������{|����
#�+b���,?���H>�`������C�0��{�%v>_)��H*D��ssD1�q-|��-�W��$~-7��K�ԈÃU�	���7��@�h�>�N�IU��3\r�-?6]_��:NϚ����vK���2O�b��B:.1��J*@��O#~�dnG�H6��T�l��[��<S*��>���e�p�^�!�-�l؎�ܴM���r�����@V*��rt�֝x�_���j�	�m�w1*z9E�e�3�~o>����]8s�vZ@��R��E��f��ڂ4����H�#��z�sJ�Lh�b g�� �8�����
�2]V�c-�0�,Ʃk!�hr�/�$Oe:B�"��G���~}����Pm
�65�vF�f�5`_h��Qcc��p�p�ٓ�f[��Rhj&��_���,t���?��b->�Ǻ$�t.�����xr�Mh##�de�d6���h-�C���t^��F�%ܒ���w��J��^����g�ɬ"8=���u8���e�3�a C�mټ�E�cԢ�g��1�\��򐧃�}�ٝ��}�{�7ށt�}���R����W���&�Z: ���p��T�	];��k�X/�%����$L4�6�	��mn��@ͣ|�0�z���;a.�&���RX��>n��;��'����{�>n�{:J�U���W��;ʃgZ.)N�(���q��u��;����B=L���p��m����cU�I��8����� ��[����ĆpV���g%�������1<�_͵�yE�u����^Ҡ�Ĥe^���'&	�G�$����YfF铒j��),(=�QkZ�>~��4.t�klw �q ,ͥ�@
} �7�6K15��7��yz�5_7�jw�k����:�[�@��gA,�o�$:��n��hr��z+i&L�!)�I�§�*ɀ��%��ttD�ק��l>��G�:;c��]ū������м"#��o�f���kK]�/�q�i�٭�ב]��Un���t����� ��pئSX�����,+���������uj�a�&t�]_K>+χ��Y�U��UrO��j>��+��CCa=8����������ţB��8�5&uE��1W���:�T����#~l��mQ��dQ�����ę����j��p&�7;ܟi�Χ��V(K0��|��=��wD���E�i�Z5�2�T�V `Z�]�3K
�ѵ�.�e�LlT)�ݹM<3�sq��_��R~�?M?�g�`3̓a^�rP��,:� 2�0[�49��C�d�����.���94��=�8�쓹=��T��F��q���:���F�	Z�%eL�L�r����	��U�� ��w�R�~�St��f�)'9<�0􎵺�I'AW��B�0`�n)��\��b��㞴@��7)� :�)�7�� �eH!���*�[@=yy��j�Y� ��k߯ ���� i�s!���#}����.L��i��SF���Fjv�G�0`�Dl��>6����/���Ub�.ˆ�X���a��"��݈�D�)���#��Feا9�+PD��U�"I�+�^�-��!W�3�b60�Cq������,	x�3��^���)����Xi�G~�Ɂ�m�q[��U5�2���vv8u9�$�L*���- O�$k��0f�I�D��*���x�E���l%�<�>G�"0ٞ1�bR�Ny�KT�/u&͐M�08��l�qj��|T��#�s˜.l�4-�<�k�X����؛�z�ڷ���LM���G��YJ\�e���E�/����v`��4U�N�X�/a8�0=!�
v�����r.�<�uT߾�-
�h�=爻�V���9��*1�#�!��攪#��u�"k(����ܼ'$���_�.]���08i�QŘ��/�T���~��1;���1��,8�gk+-c�U`�̇()����u1��R�3�����Жu(�1+��͎;�������	�1�ffg�H�г��#v��N�
���ES���*���� �` ;��`h������!-p��a�#Ȩ�#I¥�Jl]叙�3����}�B8�>&��<��^ZNMF~�P�9H��i��a�4���4J�d����m�� B�)~�΄��=_u;����I���9����ÿ[tx�l�� ���K�#�>0�a�{nV�❗m��*D_Ĳ����d�I�_�'f^�Ǟ�Д�L1���Y�jWT�0a��Yl��w'A��鿄I�w��$q��$�S��»���dPaɼ!����o�hKk���9�gc�d�~�Q��F"�}#�9��w~��Wo.�E��M��嵽ٽ����<9��s�r,�P�4�:��8ʤ�	Q�pa5�.����@.��[���87�@�f�=���l	r��ʜQ�<vdl�~�e1�3�<�
�g��V*�_���8��ҙ�4�x��*kg�^�ɓ�p�[�z$}�'b?�h ڙ4�1�~Z��3B=Z��D^����\�=�t�R
0R�=4�Mg#����&J��&=ϭRL�4VߖV�MQn<T�ſj�z+��N}��k��e��E�\����w�an��h�]@XaB7�T����G��ı^�P;dH9Fˑ�yhgS<w�b�b�Ҹ������q*�X=rrڂ����Ş�V���Vv�W^��� Z}�->�K�ꌴ��R{�	*�TI.S�X�
8!sS��?S[z�"}�I*�W�lA^�Mb�S>k?$r�k|�m }�-���Թ�p����-TJٰ���:��%�Oҋ5�`�__Y�2R���Cё�'�;�1!M�� A|� cc���0����!i3�8 }���޵��N����ָU��؃�g��?���N+T�R���܃��9�Q�#��8���؞C���Ҝ	F0�r�u�Ϸ�9	!N���e���.���@�-V�̨����q��H^p%���n\�n7�l����B!j�\�۲��a0�0������. L���o+���{y
���f0�=�NꌈAI�!�0�J�4qc�I�(����	>�*k���{�ҋ�B�*xơ�Hn��V�so֟��QDi��c���"@pV�]���lr�ΐ���)�����!M$��V���&U�SM\���|0=�����ď�PB�^�GP��������y�2��Za�������K^~�!���@2fj�1N�V��5;�7��L^g5�=����q����	[�
��:���i6C&�YlǺ��cԝ�@}��5mQ�;v�?$��B��A��w_�'�|iEk���gD@p�@��钱B�Q8N�&���K�.���&�����w��\#�[�A|?��ӗ�v,F�\�ڷ���@?Vd(D�� $}b���}M�++�Uk�{3����&��Hf�r�C�A�gL�8�_G��i|z+K��hxgsG�;[n���xJ�](T��A�M�ar~��V�=Ɍ�M�Fj"�0ǟW@d�:�o{�vZ�J�V�����ܓ���+�Vd	C<&TN�G���eo��:����{[<�]7+��ثt[�K"g8��mL��^�\[n^&���j��KI�xm�\���'�✶D�qk*Pe���ձk�g@>a��M�NAd-��j���L��L�i��n��/�2�	�����PQ�6P�� ��4���1�y`��t:�Y$��N��I��~I�`늜�^>��v��W�"��69��?�"1���\
����V���C`t"Rp)��K'�� LG?�t�l��1����rdjE>/a��a���*R�j-��\��JJ�38Mv���gJ�%HA�FUY���C��e�k"����� ��)� c��Xw�TG�O�Օ�9�!_�*QQ��M5��\$k�ɰ�;N^z�ȁ	�1�{�d��
�=��$(="�(�h\Y� 2�뒧}�X^�6�dS�#EDݓ9s��Z*���rR ��JH]�#A�~��_�N��@�l	GC�̀�E!�b%s[�+]pC���H���6I"���fy��<��ͨn�G�)=��L�wc���z�=h�E��*�N�(�A۪���������w��r��Җd�m�  �#���YO��@2 N��'�o�}��/�D����
ݷ��� Z0<֤��_'��9%�i�Ӆ��&M4�O�b7�; �|�T�JȄ��C��m��}�0���9�fɧϮ� Ԍ������2��ɾ� �ߓW%��,����^���Sk�<+��,��LÉx¶��V4�i!}*Ǉ^~!��Y��GFv[5[�hHbJ��J���]��&v�uf�&�@U���tHVL��gٜ�J�,Ї�[�=}P��-����Ε}�G���C�o�W��6�����Aě2�>\7�8�z /����	�N���DUA��Pa�[��6��?��Ō�w'ˠ��Ϧ�MoA���b��
&����hN29���Ì&H�Ye��!g�b��ǋ�8��� m#�Sgð��;#����C1�y�3z�G�M^"��̑�:1x�%���e�?�6�V�e\ʋy�$���y��
�x�p*0.��y'�J�w �"����ȩ��lD�+/N�?�3�q=�#�D�p�ɖBC��SES�
�(>���u|:��ll��Tf9����}��%Qԩ�*5���V���"��b��@�΋��|�g�$E��u��(���a��n�_KCo��P�uG�3ZE��Ae����9iDyD-�V�wI!���G�.S�qR�h>���k��H` f�L�� � ����%��ZRx��h�bR"Ä�.K�����Wa��{�8�T�^�魍�VM���2�o��E����E��6�\�Ɵ�PK:R3(}tz��U+�d@��q���iH�|�G�[�U����DJWӐ54��5q���v�ȃ"񊭒�K�P�c�A�)x�3W�*MA�*Z����p�����ldu���^�b����v��́o����J�Í$$�~[����V�ѻ(��t�)�hsb�Qp}�0@����Dkq�"�>���}A�"���ٍ5D��a�3
�quu��aIA�~�_��փ:�q�1���!U�"��v�n�[Q�ֺ�?����'��t͖i��օ��c�*J�/#��N"T��_���y��-�۷���[�:�sr�?��=�= ��Uj�!�K�x�5�iя��лF��uI)c�NbGL꽧9G�Y�^Q��?�	�ϑq)�g�*,�O��J�ɧ8��>��n����-��Y�:�	p=�ƙ�ݶ��5yO��_�ÝiW�|>�ѯ�F�J;R�W��Ge�΃�-��>'ɿ�+6U���؀~M�nK��B�k�OY+�M�~RIx.��l�$�u]�7�6�,�~��xD]��Ӓ_��Q�~�e�Id���^C&��p'4��L�9�691	Wr�E`G	�g�gT'�V�|BYC̲��^|�k�U<>Z�	Ŏy����b�tc�)e.M3gBS�D��a�92�TS��6�(Z���%�j3�B�o�a��P<�3�U�`��v��E�Z�zR)q�����q�ˌ�����6w��ir�S�0�)ډ�aS;��#n	y�+��'tį|ɍo��Sď͐A:��b�$UD7b��M�An! &�'o�꽬��Jb���*�ù�	���'�t.��C�^7}[Mz�8�� �6� h�X�U����3
��
oc�����,,���xlt�H�c�yV�c|N�e�W�:�>���('b�x��m�(£\	��os�x�6�2����-K�گ�r)S_e.q !5�96��^�#�)%MŮ=����]�L�ǔ#��A�l�p������}NHBCl	B�����ҟ���+Sw�J�n�\��!�h(�b���I����-x��8;t��S�CE��֒�p�Ԇ����3�[������Ͳ}�ӒmË]_5	Fc����sٮC���^��<w���ٻ���b���k�F��kC�P(r�t�Mf!��u+n���e�v[��0����Q�-����a�|ڮN�K98'Ło@�>��cش�똎�v��R���������I;�`t�^<���#�Ż%����p�⁋Q�-�"�5y���W\�ƽ.��H�y�$��T�t�	�?^���@Hʬ?*>�AqiS��!?=_Ir��W稕	S�[X�#��,6=@ҳ��[ڰ��&�m0緎�u���jc�D�F�c�=�GD������?9��a��D�3�.�w�ڗ�c	���c����$�Ԋ؎-�����2��G4WmyD��aZˡ~V�w��t��H̋��<�C�p�%�S�Lp��i6��B�HkX6����*,�)�dAΞz�������#;f�����=6�0�<���$fi^���'���`�j�`٤���6��8�|��@R����J��o��VՓ��u��b�J
z�ZK�.��R�g z
.Ӣm�S�NbV��' ʧf,�M8��҆gt8�I�/�"��)��A%�Z�Q �Hd�p)�_�hގ~f4_���A��8L�'9�oĎ%��R���y�����*�7�A��&u��N�W��d:���u�����~e���vO�������r��C�� ؽ��J�6T3��)�Z	
���n�˂V��g��=h�#� �x"�Q��x+�/�k�|��Bh���է	F�XIC6nasOV�� ��[wۉ���X=��#j���і�>G���M�)���\��g8�V��ۭ� ��3���Ye�fkQZ�h���ٺ	��G�����X�%x�mH:�X#�r6v-3{�0�dcs��$18旲��yH��)����[hIf~�x��ܑH4c-��.Y�����=�t���y��;o���\�]��ǻst��
���6�������e�_o�_7�a���
5�(��>�U��'f��t������+C7SSfvW��3�ƞ������w�g Ǳ4�iV7��:tWd��s\I
�hk�y��jb�y#�A����I?5��u����'���}0�S�?�g�5a�J
�A�݁U�����by��R�,�3'pH�#~iT�rSR�0�ʁU�~��)Y���%�/-g�@Mc���ǃGmQ@�)�D�}{��V����B��-��9��1y;�U�	�ͣ�w��t7��n��TNy�{���c���eS�]G���~��џQc����X���-���3%���+�H�+�"iF�G��}I��C^_�&�μ����e]�_���o��ӳ>��bd.IC��<�8�@(�QAm���x�����N�TA���8����8B$vDU��������Y+��ԮE׳�OU��-;�S��48��G\9񄭾�ׅd-�ٞt����W����#XL�Fy>�g�����QY
�FD�a�V7�40&�=J�;q��&)��A=�̫���"����fe�p��Z ��p#	In�����B+���g��0ˡB��;�(��ҿ�-p]�Q���d���G�)���G��ǚ��E��\Ϛ��i��WQ�*�~�(Gv���ǂV:��"�D��e�l�J�w;��t��R���Q�=�Ḇ�s���w|��{H~#��;c5J���
�	� �X���Gu�%�p�59��(QZ�x����QO)׸�z�/����C6ԥ�kz�C-���Q�P��49���ת��Y��NQ2��IOtQ��|e�v)����⬫Wψ�cn ��|5���#�����y���oŢc�G�*����gf>�2c�'�B��zv5�6�7�3�l�����<�����	j|w�n��zO�5���ۍ��mK8xP���ݷ��O-�<V�L2f~ǳ`�o0y(�Qf�ջ��o:��	r��Κ��xG��������4Z;�E��T�J
̝�d�U!�����	���!�?Ti|1LUp���U�3b\S��u?���~QUC(�V˛f6����C�%k[���GJ٧�CA!�*f#��X���쐢�¡��h̛�@�9WZ�J��rt�{���aT�OΠ����~N��x�Gp�1�h���Xn���\���W�\T��s���Ʒ�+��N�����B����_�hD�8]�����y�u,g�Ȇ���֋$$}��e�-��)2B�oS��6�
��ҕ^�����Y"�����K��Ǩ�h�������������pQ�l��yF
�����_�M��G�7S�sx�Y ��e�֓[��a6HT�����G���j��*�\A�w�6�҆/�̩҂�V�ތ=�IE�k�~ƪ�RO�����Ѹ�T�.������XtQ����������W�$��p{�p]K�b��[W��YL�&n��5�xлSԎB���g�9�
*w�-xHv�Y�����:E��*��������H^u9G�+�#f�����B�� f\�~��sE�/�Yߖ1\Hj���D="� ���9��ÿ�O�Z��}M)�-�NFq�O!�L��b%p����kc�o���R��p��U���|P�>��*��,���k�fW��]O���e\��������
����zI�Q䊭X��[3�u��Y���]�˕�x�[������Ozs_�$��XZ}�[��=�'P
y�~���#%�	q.���g[�ɤ<��M��5�7��Pqr��BA��D�:��D��a㺉�rK���`�7��j�wnN�u��zO���bOB��/�p�!lP���ϒ���Ǖ�U�QƤ�K-�o{�A(��#��� ���E@[9��<��|3z
l�c;*n�|��r��;�p��[$��ϜE�CFŁ�Z&�0g)��0��� <0qojDV�R�G �N���ӡ��6=�x�W��8S�J���0{>�}�(��Nd0�(�3y�%���H}Ti1rJ�N�г����&�|�	s�����I��Q+��u�3�:�96����~M�#K��}�i�!�e�6k[�]�\2S;���߅���S���d��.��n%�1��W��_���H��xi!���3�4Y�EJ8��*ӽ${����y&|&9�7������5��� �4����H�"U�H�= YB�@����3�,��Zs%K��1yO�+�?#C��D����}���W�����;	���8]��2��\b���I
�r�hQ:X�Ř'��I�x��Ȧ�#6���h��G�|��?�h�5�w9�J�FN @���9F-��"��fMx�Pm�P/0� u��+ʚ�2�z.6/U!�w�m�BV�)�g��=�h��^
V[	��L�Nd�n_������q8�#�0+�#���������r��	)�j������}c�k�񵺌�9�+-Ѽ�w�t�#�D�D?�c?��_�!����&���+�s�����J��ң?8����'>�O!�h�h��s��7��ѝ{�E� wO�q}�����;G"���6u{Đ�����A��C��Ǎׯ���_['�pQ6ߎ�� Y"��c�g��У�S}�k�'��;;�w��rQ��YM��?��3���>�r� Swf�jXl q�b�Da���5�v�����qxuqt�
vPOMJ���</Mf$Q���~�3^\��,��[ՠPf~���Xe�"�۱4�P*w�.�$�63p&�B�wʂg]M�f?a̞i�>�'ӷ �`i80�Jc�C���2�-M���gPq�^��+�kRz�o/���˅�=V��'Vw�=��%��c��کYP�wr�M�@��ܟ��6�B!�Xہ��a���R�՟@�b�9"���G�s:O�׺�<�iDj�W�3�-kS���7�}��,�� ]/�Æ�xCҴD����%ܷ¡��Y�0�5��vFj���M�6U���F�!#�b��yYR����É���U�}���sq���ӛ��[ S�c�3Tۊ�ƿ��l�6�,��R�͜o���sm�����>��;�M������a���0�d�X::n��W�W�l�S��Vu<;RlwFu�v9�HФ'�d'W�o�ŭ�U�K����}R�~�}6���׼/�e|6N5�7Ƌ&`p��V_�ꕸ���ha#��5�c7�Η �dA�v����i畛��`���1^L�G�74��w"mjW�:����1\N�r��Wڤ�|�r����2�:�=`R�~~�ѤTT�H��
����$��j�'ƍ��x�_(*X��y����}��[��,�����P��G�:�r�0�a�3T��{��B��%�(&X8��P��sE��u�;P��	�rZ����{&�'��f��89J�՞�o�Ľ�F���p��E'�_(ߗl�d-��`���ǮK5��=��V�5�V�d��O+�CI7¹!W��!��J��s�ed�~3Ns9q�Eݞ[-Hw�A܂��a2����G��+�
�:/8 ��3�׆l�T�R�_K�x�}�[K�P��l?���S�c�aQ>��adO��0�k����n����^�P%nHL���F/582O�� )�Ӄ�˧�U%�+0%ޖ��L�f^8CT� ^�^���U��p�tx����0R�zD1�,Z�o�eb����[�����fE���x\��R���������2�h��T�~]��f�
P�R7����\�WQ���5B��;��w�,a7��(:gb�Ͽ���1h���C��!} }^�^�pp��_wT���=Y<�Wze����!��:�}�<e�L���xw����58��Ϣ��Bp)�I�����;��NaT�������<d"��1��� �6�cKtf͝����3��Y��v�Hl/I_A��̚ ;Ea�����Q�u�fZA5ȵ����%����c��<,8旉��q.��*�䖌FΔЇ9�u(�ML�d0ZT�������j��&̑�e��rG^K��}���J|�y2ˋ��Jٔa��zI�B���N�e����Y�.5ҝ-���z�-O���ԍ5�M��j�إ+�����[kl'�iy2m+��V��T�߄�d7#��d�]�uP*)��&*X�.�Ӗ�	f�cE�[���ev��`��ݤX.!?��H��wZ�����N���Y#�=�P�=����hFi^N��y���^;�We��S�h��F�0���0J-�Y�-V�̐������k��w(QGJ���8@4#ϳ	Ȥx���Xp��s`n�3��iq���L��C�
�v^ym�3w���}���Aw�ޛKX���O�jy���J�Q(����.�Vΰu���s7C�p�Ax)'��ΡS�!�R�Є%u6+bN|�U:��J���a�zFÙz�?e�ZժG�����!����w9O�P��&#[�8������Hb����������d�B���N51���O��ӕ>�zw��녳!��0L���מ`�7�\3��0�vڈ��wKG�Ә2�u�䢔�ђ�T	�>-��{��lL��1�@+.����5�~��)���0F�����ۃ����n�t����b
Ho�"��8�)V >o;���i-��USFm/�,B��j����XF]�4�F0�A՜4�@��Z���Ȅ����P�<$[�b�y�@/�K��tg:��EwwD�s	ԩ�  ;/`O��J��1�X�m��u��yi���t]&Rj�c�RЉ�9w�������=9�E���ngA!�]����!�߄��:�L�Mc@���O�U���ִQ��#w|#�����_'���$�}��ؙ/^f(����Z��g��.��|#��h�g���]r�3�9��O�B2�4n8��a�l0[/:H�D�y�6�H0��_�ƒ,�H0�0N/=�6L/iat��0-�> o��b���/nsaN��@4O�<h4���H̢�6V��ך��$�:4͜<c�+B�+Ǿ���
C���̐�0�J�{B��[^,!����7OZ���� �JV�G*ʹ�n��_��jy/3VA&*�C�U�.u*��1]ve�̗H�c��Ip�1�M\D����_�{o�\�T�˞7���L@v-��Gxn��u�����8]X�3є^8'�՛��7�r	Q��[bW��_���F���H���)t��Jn�x,ZV���|w9;����Dt�F��g�熟ӭ�X?���.a$yQX�J�(ll�|�^{�������.��F7���ld�겢7h�?�Aht��I��������昼�cu�_�r�:�s+2N; �H�6�"�JRjS�1XO=�F	��5\�٢�\�űB���xU�ӂ��#I�:d�۰��H-C�\�hǬ7���4��K�m���5P�'�L�T�ӄ�5�|�`G{�2��i��Mĉ�v�/U�;*�'h�;d��,E�J�tv2t�q�Ԋ7��|{h��/�o�=\L�O?��2~�|��^��p*ٺ�g2���\���Z���G�U}��<ɴ%���ϼ�e�[XǍcV��h5o��ag���t\����n�zܾ�2|����X�|��5V�~��Ck!QѰ#6��O 5&�&#� ʻC�0�1��-���*�!�u�pJDI���m\��ϟTҲ�F��B�|�pQI��M�ix?��&�0�׶Z�Ҏ��n�-;&����te4rH����^O�`���٬�C:&ְjQչ�������0�yr�1��8���mz��
#V}b��#�*�(�@2��)�#�������{�]��(;��B-9��y��
|���R)��&�:�B�B�H��j������jc��R����:�HC����|#�/6�S�3�Q�~�]����Q���	����*�[?�>joi����A	�,��4�; ��fB�d�>x��Dv�u�FJ))d#��.�	/.ak^�����'��?u��
�֚�����%(�H6��3An�V2'���n����C�*x�o(ZeX(�#Zf��Y��l��g_����	�)ʆ�<k����'��>Kyh�yeh8�b���(���� �l~ �^�yV5Gh<�����t�-�|Fs֖�� K4J��KPcd�׏�KD� ���.y<q�<�ph�WCx��'6hdZ��ڋ���b��ڨ����ђ�D9�ʅ��x��2��zw��AR�y�]�P!�����_M��\�~AqV��r;_�v��U�Vs���C��EP/���s3� B3�6C��I���l �cBi�|�嶠�չz��ﰜ������p0G���eF��E�-y�F;8Q�<!Y�;F`IEh���n6P��m��o-V�PiܞF�"]�h7�V1]�7i��'�		�.+������_8���й�xv��	ڝ�Ր���r�0��I?�䱐��1��I�>)�R�R9w܆�ύخ�
	>�ne|�I~n:�F�4��v�C&�觋�@�]7��h�d2%t���A��xC<#��6���k90H�N�S��h��3��нQ����(���ѮO�e^��D����D�0�� vT�yn�Y�4'"gNb/}���톿�I�_B`D$��=@a����-��B�4�#��L�	N
 � �S@g���P	����/��s�T	���hy6�wBa������Ո�!�3�Jj�*���_MN'�yRŬ-��wD]�n�����>��T1}θ������fǼ,-	���/qt>�X��TǕq'���l(���Jo����C�7>����v�ާ\]u��*׉zB�m�f'�&��7�i�fc�ާ���*B�^�2ih��k�Q�
����J�6�E��DE��h)��<-���O咰p-�ź�S�Fe_�h�uΰV�O�<��o�W0ESdA��ir��:㔧���?��w:Q�v���E��Ķa�[�5�&�� �,-��x�������pPL	�"ǠwH��%>�,XM��0���s�1D}�I���燎��_�?�7��*�y�3�Por��fk�`-�DF:�H%U^�-;�A2���T<Ys��3,�_Q�֌ �Hv�"�sp���z��aD��5
2W귖
-�e�5�>��0!Y/��t����$=��I���H��:����ߋX����D�l�fҾy<n߆[;��>>7,���n��!��Ù��ї�OU����"k���o{p�`C�f��}�G�:w��?T��-� J�F��I���sPE�G�X �/�f��K}�hʔ�L�
�^7�a�5��l�x��,7g����
���2'��,o
�AZ�7�ޏ-�ė��X�/mYSM��v>��QY*��n��Pa�����_��P:��,�$���r
�A�*���������e�T�C�~�n�<L$6��c����Jy�b����|}��w���6�w�ry����Xx*�ٙ�"/�	�Sl�u4�[M����VKrŭBͣ��_�[%�m7ݔ������+?6���tH�8��5(�12-_G�l��1�נ�<p9Ή����dyO��e�Q"F�\���1��r���C�X]�qjD1�*�:�Y'�S��c"��(����"W�5J��6�����(I1�F��jrW"s�J�յ+f��?���5 �t��A�Lh*�*�PM|���r<��f�hq��}jk牔%8��w@`]p��=�yn ���[��E�+��{$�]��ܡ�/�1Q�M��m樦�X�^�;D���fS�/��z��sй�Qs�8/��KOt�Y���@(
]_�$���v�K+�bs�d�M�3��N�G�V�ڷ	 S�ն�����ٕl�`��˂��@L��/��5�	k�4�������v{�^�8t�%�>���E�>5��mȔ�J{ydt�tu���!�P����s_R��t
�$<���Q��_��d0x����/��K`'wZF9��Z
P���E�
��GZ툿�Wa�"���˫ȿ�S/�Ъ8
�)*�[nA��YS9e� �ߧ�&�7>�t�L���q*a%[�|� �gﾴ���xh8��]D�r#���Z�@��X��T=��u��q�g��q/�u���U;jn��!�^��d@)^��D�$��d�b��=��[<�x�X]�^��C�E�z~��]J���ڳ���_BT�F�'@�Q|�K/�ʚ��7-%rb�-�A������/����}6}\Xә=�������=�\������%��;�"F�L*u<��n{ �R��CŎg������1#�N��[����Uh��c�y��X18&"��&�'�3����$��7���3DX�cu'4�}�F	��B�n�+��V��i�:��������;���6�]�nhD�Ş?����]�	2�_(�|�مVW^<*'$у+�(������ɳ�N��vP��@�o��Ѣ���S����aA����ݳ�CJ��1�ޓ�O:o>?8A�o�u�̃CJv�0x�kʣG;>�h`,��j�f�2G�g������rɪ�ʐ�wNyݓ`�R��
<���sI��F+ݷ�B�Y[bL�a�7�B[a{���JLgԌ�螃h�+�s�U��͑�W��(����%ـ�J�[�?�~�^|����@r4 @���ż��ճ��{�7�]�ңK靟ӏ������%Z��OZ$�$�R^J�s�1;�t�)�1�8ipRE���&$�W�������K���|�y��.��U�N�va������,&�Kq���BPTi��x�RD���r5��t�k��a�����q���>�Y���_�M	p�6x��M)�Տ/I�-������������_N�(��N�����V%�����w����}��S^�C�^(�Y�b숔r�SYdo�9��J����8Y;O�C��~��bG���Yy��|^����豙IK�ˉ�o��?5�����$��p\�hR���,?��qo�g�j���]������|���1�Y�r��zK6}���S�l8t}�*i�:4#�Ֆ���M�;�xL�(k��Xp��G�2�'��&f�W;���>�o�A�Y-��j���t�M�.���[�>�x�
��v��#��;>-����g���� :��}�G%��O�v�(8�1��醃=�cQ�cw-�ȌUDg}��0�m�˝���-s�RC��c<�^�a�������i��^q���'��<5��7�N\~�l�d�M�:�?�ӳjs��b��ƌU���x�3�}0�5e�LeyM�o���TcI�ؒ�f�V��e\����<�9t��sb]!4�1O̹��b�H��Fˇ��4B��8`)�������2����3&��?tXg��K�����j�	�~��v.���tfËQX��ҙF����)��r���2N�>q���Y��<�f�����k��el[�:�`[E.>�	�{j�~��:`T�KV�����,|O2H�$d@���1Tzغ�y!�M|{_!��ʽG��J@��(�q��?Sy	��F����HǩѥN��o�_�GZ� �Qr�023�.R���'3h;��q&R��t׎N&�"B:��ڨ¯[�š��i0��g��2��b$I$�\Oȵ5����T�<�J���[g�<�9����ށmŜ�� v�L�����l�w�|�GXG[�;|��y��X٥�����2$[_�oE%��Xā���\�ZHh�s�'*jѸTF!5�z?(��1�����M���jP�S>G-kvC��^�]%ҖO^C���œ�\���C/N�(����ԍ?=��o�CR���w�yN�\֟a��e�AX�lq)C�q�2��=�|n���(�$Gc�H� (���\�Pߧ���}�%���Nl�ҷ�x�p�:F��cruKE�(�)ѭP�bc~- ?�w ȣ�;��	[ބ�x1�K�َ	�1t�M�p��4�L:vvےe�3EN�5�H��\�G�������!�[�#��G��%�M\�'vg��U��M.�;)e||�k��m`���D�7��C���!5wmcϻo�c��4���s{ya�+@9ի�Fr���3�;��Q�����`���{*�u�iu�������e���+Q嵲+Y����6��T��7'
!�R�2@�pI�}�7kP�e	��
�,�V�r?�m7��<i�M�@���Q��� |H Hȏ��ι�j�+��F�ÿ����*��?|�S(t���藚�w�o1L�3�ҡ�͇�Ӥ�2�t-7Ͻ}�<c;>�N��u����@��LoO����Ղ��S0C�]�G���5��d���:�H�����4��_giD�솙th��6����y�P�Tbu�*�9v��UC��7�Cr��,��9j��y��� �w}W��qH.�8GC(��է7��S��f�'�k����wd�a�TbfM���'Y�ٔʋ�,cs�g�4ـV�G^u��Y&Ȱp/f���$"\��$��%z_-�c��^2�`���9��okF ���J/n����B=m^O>�Ahy�+�"W�^�@x��0���^U�B��nzc�޾~�o�+YƓ���XWK�|����¤U�➝B0B='a�'`�%A��Qz���i������,���6�d�/�d�/����z~�Gn�wGM��f���.��$��-l/$�S	�9�JV3�o�'M�����P�o"i1p�/�R�ܮ[�P%��:K�j��s����:�4G~sэbEwH#b�Y��߁��(){��T�����9(�q��>W�~���	qo����I$��k��jG*6��e	�o�:�-�-BZ����`
|�[�E;�̕�����Dfi#�K`�i�uTu`�R�)�=�/��)jaa��l�O=8t��8����Mla�|�8���t
��1")��Y5\�U�H�+�^m����w�DH����v(�]�L��f�9�lx�������9*��L^	�uH#h�{����p��+�W;��8��}�B���q0�+s=ȶ]�շq�Nf��(��Ty�n� �tp9s���)2���2�
����9>kc�ի�'�b�zE�k�Ĳ�r�<�+���#�6H�;H�`�.�}e�*����b�z:1��v>5�w�5���෣�Ƀ����II���+}�[�,V~��״��?T�a�F��9BL�B ��;.md�g�YxW[0���_s��9u�)�4,�Т���V���0U��}4��8n�$�/Eͤ��56���|xσ��V���������Q�#u���@��?��6>��P��	�;��3h�������~pC��/)�w�=����ֹ���2��M�t�O�D��h�q�|8֩o��<��#ٍ��g��F�˄�g�ظ�� �y��uq�m���wa塀�/o�h>�W�3V��4I�ЋA��O�K͖f ���E�G���uZ��K�� "&�$����ѯ@�3�*���>�P�[˨t�zX�7�EG��NZ���l?�m���:H��0Kب �G�s�
�ƣ�P�ҧ��?��hs�.�����唤�:��@�T��2�6�N�!�F@��ug�3C8*���Ҹ���%���o�u���?1����t�c�*��Ӳ`���K�R����GpV(:5�����,=��ٳ}ݑ=2��^k���a͑M�nORh��q�OA$*WZ3�zæ���a�Lmܸ�6�M�ф����P�W��K�
�	i��Q5�tU��+%��G7"���q-C��x�[�(�i��vҸ@�cx����Ԣ��JQUy�Â+;�01]�3NI
���g��(���هG��-ۥ��
%%ZYZ}4V���OR�Vհ�%�i�r�IU5t}hjϭ���g�7ͺAvnp+��C]yN�[��||H�6�QBH.!��h�C3*wz5=ӡ�X��Y����C��~IG�~#�& ��.���Ŕ*	hE{y�j<[�96��Y�L��.����rYN��.�)��.H��|���r�����(&�YTV���!K�=n����c�L)�A���,�(�uW/��ja��{cԕ%�h��N?�~ߩ(i�䠱T���7���S�������lҎD<),ivz��|��Y��eE��1_������d�p힅�7lz�6�BqoeL7 A����m��']y�9�<�֨Z��`2,�tV�(v.`p@81P֥���е�^ѷ6��4�"�H��R�A��4�40�[#9{X1I Q�
�� [�U��Õ����_���I�O��y��<-l�Y�jp�xG5EB�բ����9/֞X�mW���@���D�B��q0N6�a�q�F���]�A��:���i�59A�(��hXOU�弢��t�BN�Hn�?���N�cל�~���\�0���T�r��;��r��l��'fao*�Y�R	�?��@��d�����5͛r�)F��
(��"z��s�!�a+�W����c�Z[����,!��`���:A�y!z�R�i.�^gp�����wg����ۂ��sܦ�D~G��U�P������<�#	|6ί;����)���;��H^��! ��?�bR�a����ｱ5���r�iW�8˦)ֿ�����~���x�H��k��x`ͷ�ƛ�����\2>�D���O���۝B7�1�CB����FQ�T<�y&�K��N� 10��J,%��(�TA�)A�`�+��~{�#�WR�9�b�ne�1-I�˥�G��=�E����0k�L��ŜT�@�5E��~�s���_����@)}2�>��l���ȳr��^��%�'��#���z$��4 �V~�B��jލ$鍘2�E\�+��C��E����cvY�IH������?M�,s��>�+��,z�)�A�M�3�khN(�Y�w[��{��
s�����$�C�V�(<�x��'�&�G߿*��am�C�|��X�A`�U~ꗏ��"&��9}A�r�ْLY?t��͟E(z��K�����#�Uқ�Y{��3�$��)K�$�d:�b�I�U	�S�_���b�ò�����d��y�z��X!�H5�8駬�ڏ�7a����2�q0, �~e��	i5ek�Ϥ��w��+��.9|0*��M�ں1��߰�|����8=X�uF��n%���ޑ��v_
�t�+_��?�w�nE��Z���kz�g�o�LT�}#)��S5hT
��9�MFB����4K<��j���)� /�n���Y(�
�v����"�nlF�����Zٙ�~O�=�e��ge�8`7ݏu`���ykWa� c]R��*b[�$uK>��z���·֐^��6Kg6��;8;R:�SF6�9"�4 ��9P����&���m��B\3h���S�i���l�Z���HLN%�P,F�:�|�h2��,=�
�9�C.C�6�aAG`2�������R]��Z�x��W��y�ĴDf��ۄU���tjr�r�C�?(b����rXN(��FH,F��X('c���'%u�<�&�����V�Jq�L�u/E��-��c0;D��f�!>�(������(��^
��qD�rO���ㆄzs��kv�G�	ǰ3g(j������,@���U�5��պ�HĐZF�_zl�% �������u�k,�aP�qd���^ץ��k�1AJ��D&d視��/�K1�-�(G���~>��+T�F3�ܬ$�0T0 ����0�X˔�B�~�m�hl��@�H
2&�����8	��O�~�T���p~�k���
4�̍�5!� l�@q�-����6�=1���œ�3�P��V�JKUв�]A2�����zf���Ì�q�[���^M�b(���-�ɸ��z1 ����P�1���[���/�d�g�d��`���Wxo�����oCk��ҡ�+_aV��0�'K�t�И�8�_�`�E7j`��_���`�Ȳ�.�C�^󶽊��l� ��yO`8 ~��#��fp���֒�ى�7&%4��r�@� �V�4�#� ����	U��І#}�
Օ"��������m��1�.��\��{;/���K~h(w k-Z��ɓ�j?`�=e�[��Ffq�=K�0������/#��g/��ʞy�1�h�I��Da.�.'r<GI�ܤs�jY���|��aW#W��7�l�o���>y�����W'�:���<�/+Փ�<�����^��.4��@ ��5*�ԎD�6��eB#��k���|ڌP�r��|P�SC�o�Ր�3�$Z�e�ʱY1���2�I1�G�]��IR��x��h��#k��	m�:B�0o�V3���
I``��J����xfN��JjN�P;7��q��c�d����Jg܃AL��i|�M\�w��(���	��֘�%�m��] [<��A �����q	����'����Y�\�Ϻ*1�.!�J�����J���P��
g�i����543��zP%���"7@��ҦM��n�zk�Nq`�S���
�s�=�(��
яE&�I�5 �=E�V�̌uiR�����ɂ��E9 c7��	���b.���K��.��ꪍ�ք��!��`_v�|������o��Sg:Sb�)[�9�8^U�M\�� $A�C��?ܛ�z�7sg�o/���J����#�2X ES�IKAN0O/�x�E��mS�G���t�T��ԣ��;x\�Ʉ<*W[-�7|�{�IX7Gd�g��{���#�r��<v�)�͆Q_M��v�7���F�^'F�\��iBT�J�@�V�!�MIp/���6�S��D߿u^g�=�����KD)����������.��W�b��P��l�|�[g0^�mՆ�q.����� �D�{-��b/�giu��T���%u�~��9���߀�vit�P���X+��g)3E�h5�¹-g���=��`X �.e�ptd�1��K�e���0�bZ�����т9&�� 3o6C�������X��O�/v@g��|�sd�׀�C3�h�`r��t߁�A]�6�_-r��������J6�$��>f<�w�ܠ���8��A�9Ș	Q�w�ɹ� y���=sz��z�]�[³�C�֣�K���0 �v�՗�U:Ӵ��焂�4� ��r�~Ёx�&p�'��ZB ��
2�B�|�y8^���卆��w��5/e߶������Ŵm<"a34j5��tml��<�
~s��(0"�6�5�E�ې����	Oy)i���x�_XТ5�����ԥ�64G�ح�J�A��,�Q��0jԁ�Ōs5~!00�hz�+z\j����f���*K��������o�1���!���6N�7/6���y�n���݋�\�Kj6<�Dv��B�xF���i]�5��v�M@�w>W����	_ܧ�^?U��������ީ�Kۡ&�:H~D�p��x�i�3�%xZ��78�;�Zw!w��J�U�0&�ǧyϤ0�Bi>��u�}���m�����m�=��t�̔��u{)"�w�ܪ�e 5��,Kn��^�i �5w���ߘ�rӎ ��/Z�/����>&_9�6��S��Nm��T�0?��SܴG�[�������nޠhe�so'ZP��\=�o�/��/&�p���O"��Ӿ2����.�� �fƥ�%�@Űv��H-����-�l{�iCd�\Z~C�3�s���ǎ`1ɔ�m�l!��"���0( M��hM6̪�(ߋ)��BD4�u٤p\O�fL
]�2\tc(y��XW騆s�2���l��%�*Gv�(b5�\�˯��W�Hh���y��w�r�1R~�W�KX�4<����ǭȣb����.UJ�"]Ps=��Ң;�ȅ�jv}?�[3����]��ξ����.����X��\�Y�r'Js��|��J]o~
�,��iY&r�k/�z^�E�nT{EgT��a�2G��7�w9�Զ|��%�$�]ÈLȷgᄋ�]�2��І��/�E�y��&���ՙ?��y�Ӱ��oъ�Lanz�3Y�~�z��``�M���$`_ĺ�w�9��Y��̺�����EV�ĝ�X�pGh����X$�G��ۢ�`��v�?���*���> ����(E�!���E�b������,v�u��֮�,-/�QW��IAj�6^��tL�U������7�g�Hi=��|є��*Ĉ׻w� ���z��x��;6k�E�-��;/z3@��� ��k�<Y/m����K��K��܈�n1��P\2�|��z�B�Y����v�<�Lf�]�ǫ��%q��1�K� ��h�����%/Q��-�\�* ��ӄ��?�ZfH4z�)r` �&d��!N�X���	��p �%���Ъ��?��-� ����i�f��k���u_�G�)�E�URh7T��"���v�sf��y~�eV�-5�ٖ�0�`Jb��.���6򞔩���a�o.�~�DIˤ<8�5"502lDM������5bah�=sK���t���n��4�D��`՜/���!��v�͇R�:�{j��.܌4Զ���Ԝ��;�: ��o�;2���I@\��s����{Ҙ&�]H��'�t��e٪L~�C·���~ڇt�iVNp0ׁ��S^%ي�k�>�/��@�KMu�x�����J�^z���E�*�e���~OJZUS})�����a�|� _^��c`;��Ay'k;���I�E���K��{� 	�Lq�k4-���X|,���5$�ƶ�C'x��dF���> Ӱz1/!���@�bQtC��m�~
aR؉��G�Eu4&�GKf�>���V�v�j,�4���6���3G%L��'+|�~6�Bh��u���Pe`���.1���(]�'����>tK`)cS�w��o�u��}���0���w����vy<�<�4`��^}���$�z��K*����>��;��p|��N�'�B�l:԰%���e!#1C��?���Bg�'� ^-<��X�Y�m���+YDB^f�rFX�"%����g�+,%�7C�A��1R����L�O�:�ME0 ��i�g`M�{Ն��ss��ϑX�D}o�in��Զ�r7ք�Ov3�sY��Sg��ék��1O��q�A� �0���|�עԟ��ϳ�I�|*������,_���O���Je["	�L�
�^���DST>�p)�Z1+��Ϥ�W����&��P`(gf�t�f��[�\���R��Dg�`���̞n�����z����<�V$�v��T <����SՀ�!�������i18��:Ƅ���i5�M���sR�m�g%�a��D-: �Zf�+��H�i�h%���c�>�mM��x�+�Y� ]NX�;Mf�zG=g�?��	`T���;f	?6P�6�D��y�)N�4����6_,��V�U_������iC]-9!�Ւr�$P�w����줆�m�Le�-��!-�(�n�1��B��K���Ol�Pi�I�� ��OJ}��{��y1��gߜ����0�jZ��$�x���5Z�{i�α��h� C����à��ˬ߰ �Y������q�Tɪ5�O�K����]���Wm4�X2L4U����>C�k���i���X@��3Y���>~
�'t�c�&E�^Mӿ�)��o���wޢ�{6dy���s�9��R�����4�V���{�X�J�I)��^{�*�g�e1-0�`
!E�q(Ƴ�5@LӲ?5��b�uH���mUH��0�:]g��?h=`N���m�5���0������SzAiTMa��k<��̕�/�kR���#����v�ّ�xo���֌N("�'t����,�P
9*D�2�4��:��,��g�kz��+����M�\�!�W���L�I� .��Mpf\�E����&O�QAj�O9f�[5�ԥo�zI>E{g��kƜp�,�!��C9���i��њ��o<E�8�,{�Η�(�d���x���y��=z�F:��W^N�)�(%�Ct;	��(�Gש����:r��$h��A��h������-����"]"��a���z�<΍y���'�꿲��ݬ5�D����8P���>���Jf�F���� �ZAjPk��/��Xe�)t���5n�V\XP�9$�D9]k�i�zJ��T#����� �MȔ��ձ���}nd<�G`2���1-�=ZA�Y�`�:����g�C��8
j�>z=6���P�� f�bD#�����`4h�"��}d��骝&*�QR�=%0�dS7X�N�b,�&�*�
�\r��'�#�X��1�B�Q�"�8�Ҍ��/EV��YR�g8�X�/��v}U�W7�q����� ��^p����s�s�� E]\\��n�
�n��!�W�VW^�8`���9V@��"Ҷ}�d�h��ezƛ���Nv{��UVȎ���ܵ2v�F`~@���$B�XȠ}���}�D�1��93�6��U��^&-�e�=�ST%섳�� ][���-o����X��a��H��7u�KB����X��(q��u�_f_��1[���$�I���@�Ig��%�I��5�a���ӎ��:w�k��KT���s�FR�I+���b�	�|���P��L��mv������Ү>�8�HU|��l_��S��g�����QX>W'��K���&陥3�c�[WoWK��m�k��o ~hƌ�_*���Jg}��)\�H{�D<��`ŔC��D�{`���w/K��`p6Zd�t�������1N��ybt�1�p]ұ��e������<Z���rj�4�kB���hNmqV�x�T������q��zX��{���Gġ3�	��ݸc���V��b�=��#M����7p�>e��-__��������:�� l��N�"�"�:1,��~�X˲�?qQ*�[�䟴@��<��4E($�)&
u~�L"g�(/o��Z���!�1�������$��+
&�u*v)��;|�-�Mc��~�Z�)C�i���a�9�{\0�/I�:T���՘�`�=/ozuQn��x@��( e�O�,�83�[�n/���"'�~�͹c�qת��I�x��W��h�a�OA94�(�%�x�������q>���t��0|���{��<V�I+�H��9����.H�@���k��Hmq���G�I?\'�]
\%�zw��A��;�}`TN�g�Jp�v{?���tB<�X�Ȥ���9�p;���������9)r�7�V�D���r���������e�@��v`Nz�Vx�B5��ؖxz	e=�!�ڢut	�j�Q��/�?ƻo��jN�������
���@�CS���cS�ز3/�B@3\�G1�i/ �*�|����@~���t!����j�����$�s��Q:|�1�מ�ھ ��QD!"�΢������.$t
�z�z�d�t��������?���4���bl)uWjJe��6��<�b�Ȥw�"���ȑ��G�$�e���<�P�����p�l\�����A�>@4�����>�z�H�ϛ� *��)�³"����@h6�~H�� V��e��v�j���5�g4P��a���k<�c8h4������m̞�>硇;N�u�S N�	F�o�Mb�Kf��Y�y��}��!�k�����%4b|G�綍����\Ԛ"�,����zY6,����U��w�c�����a�rC3��G.����!�l*{<�y\2Dy���~cr�P.<�x!�cR���=�e���ܘ�_T*&�$��nq�%'���MH��bӊQ��P<�ƅJ*-��P�`�Z�	��;����Vo��A:[]7Z7s��d�Kd�o�%��#��-�epC_1�(k�����|ͳ�����s�Z�c�2آc�nj��2�',Dus��̸����Hy���d�,�n�����#���G��L�/���{�5�ps&=��h:���RP�4G��z�!(����>p�ش0�8���|�HՇ�۾���P��V*d�����1 ���)��mfV\¹iv��;���Q�_á�HЄQ%��WGj�}M��U�/����'s-�K=��o����!ꖷIc���Q���詣���]��u�kQf'm�,%����0u`i/z�0iD=�B���{<�AGE+�V�@�٤ځ�G�o������]tH'<_�c-���l��	v�\�Lp��Ϥ���MSƿ#čfY΃�UgI��;���/`��^�-��M�ӎ#�g?53?<�on���m��Nŉ	�`:����^u���؞%n�񗷓:?� TE��[Bj��}�)�2��-Qo�`U�	lb]���jo��ؽui���@4Ѷ߳R���~�0{�^歸;S��Y������I�iX��ĢH⚰�x�`�.2�ڴe��Pǰ�yR�Pjf��3?X}0_*M���L�����0�)�*M�"]��mi�w�8EE�l
�B-g]'{h�u��œcQ���#}>E�m`_�_��e�Fz�?�.�{���W=:�[��3n���xg�!��Q:̧UD��L��,D�\{j\D�� ܵ��:#I�b-4����-�q#��2z��������%���޻���V�u�d�I)$[hp�K�*��$;mj�����.p@,��B�yE�ewA;`%��M�\[a�U�"Ѐ]�N�?@�l��)���ޓ��O/����!X6�$�#�ZWA�f�9jW6��?AQ!yx��}���VT
C��cB[�W��
)4���Dʃ�~1>�GE���Ѡ��I�R)DF8���b�(z(ö-OI��/RYxM���Z̋�DB�s}�qK��$)�/���e}"�@ҳ��q�%��M�z5�m��S��5aQQ��T�����J�.�d�
�V�!�����0b�p�Y�Kn�|)TsJH���(k�U��Bl�(�LWD�Q�nj��E�(|?��LTm�ܬu"X��a�3Ч�Ό� P4��	�H�<IH����h"(:�����M{~���Ht2�8�X`����-~Y>g
�}���p���=@���D u�[��K�ǧ�HT&��Ͳ�<r��.��
��4psdX����y�s��m�I_�q��')���A�/�E~��<}���8�z�t^�$�g��O��^Bz��D��&ɖX ���"��U�&�������E���&�[���_����p��� w�Y�N�Zhh�z\�;s��Z��&H=�v�� �ށ=�v�i��?sT��g�l��޷�V=|��� 9�4�x/��>bKC�����'#����vuB̩����7�`��`��F�O{����;�T��f߽ꝄI8��5E�G�W�I	���������b�>2Audo�����C��lZ� ��Z.A���o�(�j23��������*�`&c��2���O#e��� �]�^��}�˷�M���-(@��Lv
>Z$S����2Z��
c������=))��ף슊�����vy7=w��v�Ш���������
vf�V��\��ߦ��d�5�i1}��W����H�1DSn�;�F�/�E"����y�_�祦�	˪;/�?�S\����b��][��jm�����C_@�OL#�%%ɸ98lF�-I���t0z	7�5>η\�r6_��l�KJ�0bT�Z��Z.���k�j޶N��j��3�s�a��g�9lV�->{�n,4`ˏ�����@�=�"6�!��7�p�>����T��I򝀖R��:h�B��-� �ET�õ4�����C��R=�6-�9��M(��Y��6�ϼ��;+v\�W��
�=�0��yv	i��?�%+��d$��i��XQE�t���ֵ+�A�S8m�b�Z0�#�l���j4H�yb����g��Q�(�������6���p��>vb�����4Ք�,�9�b����7�ȇY�d�z2#�:"���%:�5��ᎁ�B�)~��Zoiv��<Up�Ӟsឋ|�-p�0�������Z'ĸ]]��s�#������.B� ')��C�*��ϼ�w+D��Xk�7V��n��)�.�]���V�p&�N�"!�oD��P����8l��=�=�L�w�W��D��#�A�o|J>;�I�Ҭc�cb�	��L��״�-�,3��X�{Ek}})@�x���L�;4�,�]'��tIU&�1�5�x�(W��NA%U�_9	�$'��2�	n_��|�9��
o�=TP�9���x����/�=�C�=��Y�)0 �!�}H�Cg<
>9��X^��� iuv�����Ͳ����4��2N]�>� �.;b�XK�m��~+Px9�g�M�۹f�:	�����
0
�z��mFGT.��Ĉ`������^�p7�L�߲��0�+�XΈW��D�� �yQ��f����l�|gТ^`q��|:�$z�6���FV�.S����Df\
JG�b���e1��|�`�\�>C΢��5SV�N�s��<#*�p�	^T2do���,�|��{��'b�SřmY��y^ �/F��A"�NS��J�k�|B9��	0j���E��N��1�]�Npc4Kv�t:o��0"`����|Y!����.KJ��@�l��׬�
�
�(My���_��C��<��b'�cG�������UN\�jn=��:>�wr1L�l�J0�g� {�t��B��d�$N�)�S"��+�_�wj0\�C�������mX\d)�;� �����Y
y�/\����~�+�����D��T��߷���յW�S��6~�)n�~����Ē��gW�C! v��PEy��fА��j:��3I�f`93�@�KF�^���Q �+���,�qg��b��� *�Kz�F����U�F<�(_ž�-����b�������&��@�e/b=f.*w���"Oo�����G�	�c{��+��6۾�]Z��I�Q���OmO��Ѕx�WɃm��2�׃�F��m{��`����L0��by�Z^#)��x�|��j\��$D�E;e]�:���C��<���:��?�]���U�}/]^r���_ܝ�K����?ĒTH�u�C�٧؍�T�p͕�*�kl�ט"?
�f�S�Z[�)V��l/�m,�`�C�B��U@�yZ�Z�J�o��Zk���%1M�GG�[<&��O�D.����8Θ�>�ѯ�Of��D/s�N��ש�1{��Z����C/g������X�R������rU�Qr0 mSŊ:��]�^ɝ������O�<��}`�b�����6�(��]k����m�(^6ęKN���3dT������`<GF���/����O���R�Vv�xQ�Z@�����K�_Y@(o:�sj?����$iw�M�T$�Ӑ�K?�X�q�H?Lft>��X�Ő��a�T|S����r˚�oO9�Gj�z�A>q|9h���g�E�����操���`��=L�Jd	P��B�@�~c���3�kh���4�־^j0�y��A֓�`C����칐��o	���i4��3��Z��b���2
��K��u�]�Q�N������p(EQ�9m<�U#�B�n�wn�%����0��Ih��&�$Ǵ�n�����6a���lJ�٣�auօ\wn*�E�n]$����*7��!i����sn��8�u���5ʤeQ߉�g\s��61�
����],FK�j�LvT��u�LyY+�����I�͎��JN�d"<�"������a����^����V���]�u9�R�w=+�ǁ��H�!�-n�u|�:���e�ٙr��Iˉ`<d��v����zy�@y��7�$�Z��N(��������[����<'��d�������e����f*q��Mb�ZLbzoy����wh�e,��El3��'��X�e�e� ȉ�!:冲����d�	��7l�;���~t
��C�O��|obH�`�r���v4�}�u�+�s�f�����7�\׻�q�F��X���2dU,~�*��O���ٸ�N�6�X�k�QA��-i�ȡ�E�-��*q�OKm�}ikQۈD���L�;,�v�>cҠ��Я�[H�%l`�vu3� ��m���@�� x'z���H[t)�>@cW.N�I��:�=~;�/^���pa��e��70ᕀ����m{��^��V���Rg��%���dɢ<_�P��х�M�/[H��$��$�ʡ����}u6���C��@�!.[�����%�0��U/ܪ�+�4�"[\�M�M�&%�u�py�.��G&�֙�V M��U1.VV�~((�Nj����3׈�v�M�S_O�7��&c��-PB[�J���.N��5a�qw��f+�Đ���noGS���������Ү���P�Y������J%0�#iS̕�����R���{Zm�{��*�<��������ls$��I�| 糍u>Zvm��ss�&��6�|&Cj��e�70�����p+��ɒ�5r>J�f5��?����B��"����1.���ǝ���I1�E��"����#� �@@Ҭ���B�3��/��?-��Ce�Q*���Qk=�~����h��Z���>C����o�d���HX��T\%(��@��/M�^`Z4O�2� ����u���Y�.�Nö�ic\&.��+�.t��+CA��Oy�����k��D��]�JO�����8����n��s��;�%gb:���gَf��F!S1�a�
JmK�;����6�2��i���x��5*��f�i_�ك�Y��� ��T�<�T�e!��_��(��7FCq�}����0z��*4���v�����2��U3�$�#���e���0��Jm����N�d��)��� 03[Sr �2�|ɢ���bD&���54G�K��}e��>��H�m]W9�o-����M��!�SLWx��P���Ǻs�"00�t�TPh����n�X� ��� ��(0�w�]�y>QG��څ�oŢ�JP���%3�����&U��}ȪH�/HV�������*6dpn�a��5d�e����Y5��ݟA:u�'�����0s9�:p����������ۢ�D7R0;��'���nΈzm�
���F�\_�ų�ǡ�D�u1���)pjL��x�W�La�f�@��%�x	�˲a�=��{c0p����¼��vq�"Д��2I';�y�����#��q�c��}��ֱ�&C����PP�"=��V�PZ�_��?o1��WY�X����~%�����Yɳ�#5%v��ݽ>�CI���M!�R"�2�n�N�Fi[��\��Ҧ1�ob�ʻ��+�~��&o ������T�@F�Wva�~D����^�9$.�8e�q�}w"t��|\��S ����n����Ў���Pm�AQlӒ�5� �w��� �����0�鑨�"�|��E�������rR����/���YB��(� �_�J:���f�W�=so�9|r�6 l������Ӵ��J�9�5�-t�.l/�Ug���@|�Еgz���w��Q=,FU����|�Jtr��U
Z���/E��~��İ�Uv�Z�I�*�q���؀�3��3���t�8y`�~������c�b�]8f`��\���7� @��4DL����*)G0o&��	��kD��������$����
�����}��۱Ǩ�G��2�4>ЌNV�/��E���0��n`M/������0kh�!�o��ȉ(f{wĨc�d�	l���d o����Y��L9$��ȴ�A����)��L���gaQ,,���K�Cy|�՛�6����խ*��bk��.�o&���V�L�<�B�yZ�b���f�;�U��:����.�N�]�vA����F��p�bŞ9~L��6 �h��?Ά�XT���R�ȫ3J�o�:� �	7%URR�k�v����B6a�8[|��RV�4ԨPѽPĒ��o_�ߝs,�il˅�0,fs���[C3�s�ZŐ�5����6�_�.�$�(�����GZ�Z$Dq�E�	e&���P��LF�7���$�W����+�S�O1?Mr�ɔ~��c$��'�>F�����_���oo�d`ꬷj���%��:�ֶ��Ğ���g>hV,����d�ZCY��?Y��<��v�R���"��Q�{�Ndz `�+���+�>�z^�G{gH5X��Nc��/��n"9�o�n��z�aHT��<=��Q�m&����Oç���\��y��WF�q��]�ςZ�\����"���^%�����&�/��Ah�荩�i�Z��^��w���)IM��'M��ܧ��@(O�FoBӚKo�<�:xA`��"�@�*궟���7�"
`�/A�ej�5ퟌ���a1���2���k�NA�]�?ųMAW%V��(�$��9�Nµ�~\������ws�t7~���A�ںC�F��?�x�v���43i�vw�@������+�>�dV�lX?�P$4�N���H���۠k�Gl|��?��H1>-Y!Đ���]rظ!%���%�RO2*է�*���J�1UϿ��ah�߰�'���2�\mo���(�����G@U'�o�6��~!y�If�_�LŒ��1�,�Ύp��"�Oou KVzhJ�:c����C��6S9�v����g��	m�´Gj����gJ�(�:��������\0�S�S�2!��(`�Y��������V�a�����. �I엜�Ĺ5�#橞/�*12p���@ɯ�њ+'��J�N|ޛ��cF�	�a��Z�Q��c�p�*;�_��옸�6��˜�!���ۆ����c/���m�-���E4��sni���5�dK\U
����}�)V6�Ʊ�]��������m����"Mo�3��[����?Z?�Q([Ggi@9Vm�^%P�Ć�(Z�]S� ���(��Ċup�����'.*c�.?�I�bB����3�z�����������>5�ў�Tz,�-�ͱBH�X�����s�q0s�����1�j�z�9'^�Y�M��h�!�Tƛ�7�yY���r����X���O�s��nEV0o���:ǈ4����isNjN[�ϹB:Z1C%�Ч��,?.#F�`��r"�//�� N��q��j�ҡ͜$�X���&T�¯pG�2���&�Ȯ`u|T�(cB����K�Zʠ�]��nb�>�� V�B�+P]��:�_��5`[���gpr�(��&abu�|��NS`(�D$x�p����U��_�b3��zY�+ܒ)3�潡�b%���Hľ����o,�\�O�|T�Z�e������?�������z ������UQ�D�Q0��SM�5r{���(&���kVyX�l[Ķ�k�O*����^A�htm`Š��X�.����S�ȍ� [h\��H����9�8�,VI&B����\ޚ�������?G����%�ayW#��ǩId���eؒBr*�������b,r10F�0ʐ�F��F�)"���tq'��m�@���Uo,�P}�O>��g0qү	yb=�����x�e�n�����u*�k[+I0��g���+�<�LbW�_�B7�<�/Qc:�$ې������c%�]@�z��y����^_�Cw獢�/��E�z{�Nn�¬�;�������_��7���4�;r(���>�'t\�1���q�ȶ"~3"�kg�~S�w_�c�9�[��bi�ڌ�Rσ/��n�r	ر_N{��+��"���Y'CU�@�X����,��(��W�1w���a�.��mM��z�����CXH�WM&���.^�v�+��^9}�K�KH�3��������eO%��s����˥���bZ �n�:F1�_��x�L�W�V��P6U/���"�𴙹��GUU0_f#	0��FmZհ��+�]�n�>�Fee�rn.�I,��#�Rs��Ϯ��,�e�ˉ�v��P�i�z#�Ş�����ekv_��VޮB��%����`����^6W�Ƃ�?�2G�_x��5n�J�	�X;�*��+��M>���E�?`�Ft�-p�Oz(u�zR�9�e�E������a���U\�K�
¶�?�7�z�*�zkp�X�� ��%#��4<�ގ�k_^��*K
�A|������,�=�����ejf�ȸ�[�Agyd5��/�*����(���D'A���fߔ�� �&��W�j��.�I�/���MM����3e���D���j�q��a�HX���F��9D���b�Ԗ1\7��o!�`�$��v*�8�+�I0ʰ���7�#�Ob�B�G�2��.�!<Z�Eئ�(]uj��֌8 �����J*g�����/��y���ƌ�ݸ�H9����J<q�6��1�a�����K��h�S��'�; Q��eZ�c�Uz�g��zYa���e:�YMBR� �� n��rDd��M�1/vI�Wcu��Iu?T0���kj/�Ѐ����Y�~�l�6����c8��]d����A�&�.lr��Q�Y��i���TtX?�8`^!ҙ�"5��E��>D��԰����^�Ed�ᒦ�y0or��v�K�� � ���M��afO��q���Bq� O�	�\c21z�d��a�L�#������f܀�Y�I^l�g��[��C�[A.�+3� Q�ʪiV�`l��{��I7�Y�͹���.80QH=�k[�2$Gm�r����r������9�/%඼��A��-��؀ͱ,\M�|X��q�#�����O�;�!1��̝֕��J[��������y����,���l�zV&�Iu�M����Z�n��,)��J&O���1v25&�K�M ���K�	b���I�Z+�;z8�}>�ɔ��V��(ړ���# �n%'�d4�F�l���M�_��j���9����Z���Y���׮�5O(�T����:5���/���8%���y.}Ȯ�x$q��)xw>�!˸�L*2�{��&3�'�����Lh�y�y�RcW�h
b�Z\~iO]�z�N���ߕZ}����)<I�q�ךO�
ó5#7���q���r_$a9��/!�@Q��N�]��|݃# t_C��0�����G*�Ԑ�����ݷL���?gS�����2^>���1s����j��"rPa��x��zx�׃?�%��6���������N��Z ����қP����9P�����'�7n�S���{0�I�i�-��a����%�B
���t��e��ɗk�殞�M�!�.lE�H֠S��{4!�3j��}��S��E~�5ݶ��~�;�m������VŃ6�sԢj�w����ܚl��5�HG)�BE�64�.4�s�I���1bA�������a@��7K�k��}]m=-tc"~��T�BJ��G窣EY��:��l�C�p��5Ц�|�����_��~}V��Y�Q���>�\x�C�I�e�`T���bn����<�v��Ÿ���Y� -�N���<�漛���]�T�Z:v��a?x�ck�����LK�؄!?8���e�>zk�q:���zw�$[��	|	k�[�{N룸^Te�9	�]sV���_:Ӆ��H��xÇ�|=�1.;��vPދ�K�3� ��E�VS7<�����w�x�@'�3z�����Q��(���`��g�y��R�9�>[G��g�����w�8��*}cu4g�o������qu�H��`9�[�C�Qz�}�֒r��m�G?�BՌ����m'��	�_mFqxx����J�u�u ]����o�������Q9?��*ޖ�kch3�]`SC��2�#�6ͯx���B_���Ҳ�|B���a�Ԑ��\�`�"?$ ^�R�K-9��'b��<��F���л��r���koA���M]������7���>G�l��A���gVqʏ�N��ȡ8D챆֙��M.["×�75��L+�Sm�f�1z�H9�h~��v�:פ0|������� �P�B3MX�F�ԲKڧ$�cfm^��v���C� 䁤�/(�Հ�T{	���#�;py�RV��?{��tI�
�[�Il&+t�Z��g����V�䝃~�/m�V�qP�!�Z���M�z�/~�!�0zG�T!V���|o`�H�G=q�K��Rbe֡?#s ��1�Į_�n�h�E �ֶ�TG�]H�>>�U��ϖ���5��i�	�D/@SI������.���x��%�T�ç\��09.vI��f�Eq�O�� ����^�~d.����Z�u7��nּ�ÿ�ڝ�L�/8ׂ��ݞ	�H�U�J�V�%�W�.�[��A$�]�{N����:\YnsB'�Ux��k^�i ��Hg�z�k�;^�����{Z��4��-J��ZL��ھ�gPֺO�8�p���y[�t�j*v@ma£x�����M��a��
��y0�Α�A���-�V��GC�T��s%?���e0����s�Z#k�+�y �Y �%����j\k#�K�8k����Gb��+�<�G���B�>ap��fe�-���X�o�5J\[����,���i}����<�"Y)ޘ@|F#�7 t��rˡ�X���/jݜ��PY��J��1uB�{}{I�VkrDM��z�B��5�;�o�b˞ց��p��B���2��y������R�}��ʁ��{�4r����G���m��:�9�n)�;����i�l��G�
yTy/�O�y�kK�<��V�@J��C̒+V�~�B�M6	��F���KY��Cd_��o��3�����X-�_�1�hr3�p�	Yv��n�~�9����݌-a���ZIxt&v��09����1qK��}8 Ś���iA�ℼ&�`'k�T�
�q��	s���-������l�c#�<Vd3�Qa}�!tפ^f��.ӬfFQ:V�A��v��1����C�E�°�<��w5�<���K<*#���.�t�75P�,E˱DIN�e���u��M?��#ߘ��.e�,���[��PQ�Q-�fo���u��m�X �:����Ø���
/K;�&J��[�c�\���>X�5f*V�;V-������װy�B}_r��*#؉��v���^���!wȺ� ���aq��w���׈�[�;WN��L�V?oش�����B��M�B�vh��"��p�~����)BͬL|W�R)��W9�Jk�U"�,�/T��2]�\�n�����P�)g�K�XB8�:N�6�D�[`��	m5���#�@�%�_Q���!d�M����#�EV;�c����gK��q2t͌����6@�zv�
<%v�QB���� �穟�s�-��ؗߌc��TcQ�8.US��ˆ�3�C�GZ�wD��311T#������:���P��DuѸ� �m�D�z�!wd���SM,���M���9����
K��� ���7�U� �-h�Kݑ�_hIЗ���`������X�D~�����6�C�ڷt"��V��ً�&0�%^m�����,T	�{E�*	b�p�f���,Α���ӽ�+7�����V�x�d�TV�5���z_�����A�?x)�v�QS�T���b�VX����-��@~D[���#M]����hX��oLP��Oy5^�`~�M�y�����Y���j+��N;a�A�!�ބ����bԉ:k�Ҋ#S�Z��Lo�����l��-/����X՗߫Q��B���;^����<s"N1\��ȵw�?6�9���RCw��ᒚ��U�'�BL����v��|�l�3���C����A���6��A��~b[�K�p��y �s���W,�kD�D�Sj�4��l _B��b� �̏���R���&��u^�X�W&��9ɏ�;El79�e��3E�c��z���闣P&��Z���U5��<?��	W��/~T^z��-$A
�����QB����E/q�G2|:QFw�dO���<�����,a��U�t���Υl�9�3b�O�o�z����1:�@�P����$�1Wݎـa��7 �;���}������^�i '��g��~-� �2q���6Jt�/Jx��W�Vͦ���x��?x�#E�g5<��D����x��إ6���n�Zf�8��Ʀ6X#w�`�VT���5 � �Z�[m�z�u�<�㙀{�;�q�"¦x����1~T�uW�?���؜.� ��*��F!KJ����\�dc�2�����g�C�}���
�v�h({g���h�4�õ�#���G��J2�A���{s2�]{Q,�X	Dxe���FB7�;?���\M t,�<4���e|_�`�׾�
ٳ�5�F]ޗ1�Ԣ(ܓw��ܽ��ѱ�gG��b_+��/GA$ %z�̈�.�K +�T�M��vS���Qj��
<H�6��/���b�c�Zm���Ή��m�&�dC���-Ŏ�IC�����G^[��9Rw!.��M�-�4{��ǔ9�c�VM6(m:�O�힒�7���_O�s��Hg+G| ��;r�@D��QN��N�YS��=�T���3ڼ��a�N� �U�R��L�܂�(^$v��I��~^�>���x=�NEO*J���7��f�����O��yֵ�ϊ�R�A�<�:�p �ʙ�^�=rY���N�f�_���%�j`^t��N!���ͫ�K*�.�ȼ3)�<N���`� H�n#�W���S�����Yk�П���Z�!$&w.ǋ���8�r6��".���(�'8�4��D�^g�-�U?����&���\��G�-��%�y���#0tg���,Z/[�}T�e�M@~�~z��(vY���0�e����L�;��2ඣ�D�"�u�|�TuD���Z��)�i�d�^i�:�+ڔ�ʂI��D�ؐ�i߿h.���r6֥�p������@��^���T3�v����f8Y��t�ߠ/tB'=����Fr�pn�G����i�go�v���/��#(L����� ���s&gJ;H+R-��i�
kԕ�J7n��\�*A�/�9�,.A*�
�vCڷ
��8��O�[�7�矕2h)��3"�m�i�Eg3��Ë��$|�P<�H�O�S ��ng���3��th�;�.����4e�ݣ[�3������5���0�G�%��HOD@�\z^��$'����)-��cZ�a6*j�E!��OC�k��>�F�A�r���a�^�@��G�qsI����b���Xⅺ���M�����"�-+#��u����S��c�?���~GX�4_/;�����/o�<a���*+M\����s��v��˃^s�M� �;I��)7{�Aq���Q�P/�;�� �x쳕�"JsOv�
�+��@g��i�BZ[�mT��fD���-1 �D��CP9<z/1G�s�}k]�PQ�m6����|��������$8M�k�������$<*w[�K��~�׍P�_�@�JMy� }��xT�ؖ���ɘ�ki
��:[hμ�eϴ��� L+�J[���*��.�>�`G�WW<�&�JsY�hӽx}�'��4Yt�2˳m��Sg\�?؁1���7h\e�����#fN�w� ��&WHB*��1�0�W��������d�X��b��l�����7�8)�Sa����I��*�M�y|�7�>z�^Nb���l�٭4�]�npR�j����j��f�h=�&E����;'vX�>����M����[�JX~_��	��N=bg�^1�	�e������*Ii&_S�h$�p�z4�����!�@���)P������gU����U΍�I��+�N����Hûmv@�Υy�p_��䴆d$K�h�X\#�t�\�?L��\�O�@_��D�SX�c�}w��RS��8���"Ug���0f:��g՟l�0�c5������c�'&�7VotUj-�^�A�0��
pS!}}�����հ�����.h�U"+����x��J&!�
�����jn0/Xd�͵>��2�a��5��~�<�hǱj�O��L������o�IBpo�^�u]���o�g��㞒ѿ�8y����T�1\��(I������0vJ��7�h��^��2�&
6������ok�|s�����HZ���tY�2oh}��e�Hc�1�l�c���#��zP�	���<�{����I؏j����B��׌:�p1�A��d�iU���.�f�n���[h�H�U�ʝq5<��.	�x��6b0�[�Vԝ*�ulfs�3���ڠ��;�w����?vX_n�G`�p�A1'���v�ԙ%s�ٸ�) �bq�p�F��/�R�%\4�Ci�I��E���P� [7�3f�U���(kGr�8��a��ii�%_A�}���_#>����E6]��!�|�����@��� .�,
�F�U�A�����\m[j��|�t���PP��R�����_ic�]�Y,J���/�.Q|���P<�8>I�3�'3�%��I�[x�����w�� �~��jY��%����s/��或Ж�'1������C��b�J3R�I̎/]��P'Z2�����)2
�4G?�b�Q��]�
.�±���;(��"�VF�D�J�'�n	Ros�"
7�8.��ð�Smj��[b;��R#��J·��^d�P�1([��^s��٤��+��ߴx����WPPup	�)�(�������l�36T�{#ՠ��r���ۙ��A92m'���ԚS��x-�2^��k���t���t���s�m�C��}I�KC Xː�hㅵ<��2T�Um�cZp]PH���	׷��ƅ��z�G�µ�~Wȋ�?��+Y�h�R:j��Ttբw\#�w��� ���!�8g~]YG ����}�  /NG�]��Σ�*EFa��8���[6B	lQ9��WB1p@��.Y�[�$����
r�o'h���r�zp�n��T�����Mi��2zGk$������'�[U�d/��~���n����w(a�v0�L�h)[w�n�kJ0�͒8j�ו�� � /�oW)UJzK�KS��%!�6�SVg+��.�F^Q)}]ad���A`��]�C!1�k�8��x���űS)�#h�Y� ��fĨ��N6���>�]֊wlL�A�-'����~J��6�r	ᄅ	S�ue�A�#f�m;YS5ۺҵb��.Fh�ѹ6ӭ0h�m��_�o��=3BT�H,�����\�B�}�����)�q(�6d��&|��9�������q�����JN�Cת��xB�����;�L��ZDAk�
x��]te1�?�P{���v(O�����U��E��3��)%�=�I�u!�?I`\�J&&}�KX��w`ay��̲%�xu��ș7�bX�A;k�C�~R���bӀ�<��������0GYX�a}�j3��:�o��QyQ�]B6�v�N+�`���zI��ݦ��I��D<�������	��U��]e��.���G�M�H�5+6p�Y�[���t��,z��o
u9�.7���6�Z���Q� tAVdF~D���Q�Wϝ�q&u�6�H��A�#I2�fȌ$SD$���R��S��:*n���������X] 0�ۈۦ�%աt�Y��|�� w��Bqe�i��?�a��{.�('�SbP�-gM&��uBB����.��toT��J��U���Fg���l	��؋�Zu�Ȉ��`=DM�#��U��N7�gp�'�R̈�H@l�<?����)R� �<��Ca�;f��R�Q��X@�X#�=`C"��p.�KT��ɸ���@z>�B%�Y95Lԏ߯�<�2��1�Ւ��95��ö������]k����� ]0��Y��tm����,�I�T܈1�1CfZ	�>�����m�=��C��dj^��ެ1#����k�Jy+�ȼt���z'��P������s3��3=u�G��S�~B��cx���yȍ�S�	]~h!�b?v�A�nlؤ�'��XG�q�$���h�(��=���B���p-~�_?���>ڎ�騄[LX+���oE����!�I�M�	4����� �r�5���}��!��0��?nyMկN�L���-�ԉX8��@K�,3���ՆD	c��w��޴� \#�܃������o� ��t��ŰR�����=(���|6����k��5�����R�Ts��a>�:>�,%z��7�
Wvĕ��]={s3~}Z�$�':���@��y:�H��^�ZZ���շ�ai�z�,���7�-�#�<�̥
�ʟ�O�P�-n�G��)V�%�@��?jR�Z�s��{7�ʨ�ƥhC�z.�E���r5<δ��9�yQ�j"l6Gi�$9�f8�N�p���[�4�Ɨ"�_ $��5�\��>Q�m���Ʀ2�$��z�Tٽ���z��O f�m�n��qfp͍Ձ����4�f�ڜ�v��\Y �NZLe�<�hqWZ�b��x#�*�E���]�%��d�!�7kZ��ֵϴ��E�ھ�*Q��A�6��J4�/=��5>U@S��Y�<������Hgi3D�=�Q�=A�H����Wg���7�.����I��i�kA��5���6cEm�!�2ߙ�L�"�X�NL`B�<qF�;���([$uE>5���F��&�@���e][ ��gL�'i��	LZ>LZ7��`�-M&Ynk[�5��HI��G��S%��r�V����V�̖�0Vj>��^�͌c����xzW971�	�Ͼ8MT��huf���S�X�ielDvxٳ��NL���N[����b��7���-�%�eto~ۈ-�6�_)��M��D|RS���ޅQ�e��=[ʧc�*�q=k��G�Uj|�E���@���R�ڜ��6u����A����*���E<��4�Yn��wcp#\�y�׃�$d��S߽!>��C�<w2��Q��U4}���!B�d�Du���.!5��.�Q62HU�1���ѹ|D�t�jq'A�R�$���~�z F<��M����e�D寧�>�J�#?���MS��5-�!�M��a[1��~� �CH٢���6:�q�T�X+�����9���&�$ax�6�v�m��<E�v��G�3̮HxJ�����«�9��Z:Bt�`�~E�|12�t�]l�!<8�+0�i,�Է.� :++�"�υ�S?��͜� �?��HL7�FT��lY�R*%�������IG��\�� b�t�r,�jj��k����e"�cTO�E��'[L�(��<�	���]��Җ)^^OJt
%�'��>�#�I�?�g9*�_�s7�ț�<�oMHU�">7:�+B��Iu�e�f��EB\B�~h"^��D.w�P��in��p�N��,>IK���zl�a��զ��PY�I0���j^�f��H�ز�����?bW� ��t�rW'�d\'��p���<�t�0���:�;��g��;��Z�2lށ�e�Ȑ�����Kw$#�r �����fA���sM9���%zcf2��H�E��p�i�\��MWiA}n��<L%!���g1iI����_�N0���k-l�76R�1�Z��{�ˈ}~�P+$|��}hlF���-T��<�j�״�=3�I5�=�)4(YqL�M@�aa�kPO׬��gIBm���ϊ=���6KNkvSF8	�������4͓^mopk�o�����[�m�XF]��������A\"����˃�\������/ъK�h<N�����}��t�\;� {z��X :���7\�+�d�˸��-�a���R�z��K_��nD��q�I��_d�����X�c���EvTr�%_mt�d�������y����Pf�6��Pm��jd��4�69Se4w�,�Aq�1�Z�����/Y���C����ظ�8�|�;�H)��!s�U�#1檜W�N6C�Poq���N�h��4CF�۪stW9�)���F��cz��3J�'z�k�sʾ�&� pd�2:�NW>��vct��|v~'r3�Ð��M�POq!���� ݞw,�]H��`���͓^��@=���j�^*-֞/�qmV,��Xf�uT-���m���g<�Q4�&�n�A�jɨn����̧͖Cπ4�N*c�F!j�D�j|�ofV�d�h�:�JN�����y��
<�z�@P��7���<)�6�c^Jx�����%�8[�NI&xy����z��P|g�s�.�L�=}�x�X��U��y<�8���^'C��y꼑o5�U���̵vI�ޜtc���{m�Du���jHP����F�=���Y������Q�,b��)6�y���U���Y�$�kz�jK��8wr��8����p�)=�KSQ��;k�<�Z��&��c�Js�4�R����`1�9j-�1���5��I\U &6��6c:��и�%�Z�I9dg��,6J�������Ho8���|e�O��s��^�ƚh���1zpѲC�w�U��m�PڸF�u��Ȇ�{>A$�x�nBE���~�+z���d���{Wt��Z�$d7Ig�=XY �w�c��X$欎�I)� �s� �����	a���˶�U�R���q��ù����FT��M�@��_؂!����m���џb�h`͠E����y�x��U��kj���9��p#7��Y�:�+����`��҆R��1��^Y^Iҝ_��`�}�4`zD�g|M�����	�w�����K��}�U��8
/E���~>e��&��/�X �#m���'�o�����슀�N�(��P��5B[�W8�=W��S�5s��q�e���Pٚ*-����$�"2T�X�2D�P�]���8�K�3�����*�{�����\�i(�b2Q�r�!��$`����4'd(�m@�8LXd=�x�9��ߨ�����lě-'�p�����d��/� ���oW!�T^vm#�M�U��U�T�2����J�2�ON����/��Q}⤡c�sl��KafŤwju��yk�?XE��T;�/y�2�S��K�h��p,��1[2E��^3Y	����<��,��xe �D��$n��+ӧ&0숭k���6+d�B'B�&!Ah����8����q^����&l�;i46�*�B�z7
��,�n�y'�د\�Ԋ�zLڥ�#��Ϙ�\>�UKt5��$��b�y����X����ĝ�yݜ�ڋ/g�̉�|�@i	��M��69h��3��ē`�,'��et��'��%/bз�>�R��@4< �grc�w%�먮����wB�c���<�� ���(2�?[	�	�;}�-�(y�2:�L�)�A,���R�@���x�8y$��$�[�tOv�o���Н$�X�h{����S���8���;�щA��)jĕ\��z�A'f��e�{Ê\����*d����à�1YJ�Gj�� ��s'{�[5���ζr쎕Fm���+�*F�t��w]�����tqb�C����&b�������ۈ���ߛ����D��TN�;.۱�p��;��iWc�s����̧���hYL�N��Ϯ�u�L]���t묠Μ�f�{�Wf��1Q�Ʊ�%)p��l�={�F̒�D���Yt��ƈ�V2T��p�5��� �Q�oK�b�PJu�*
(���hfy/��^�ψK�,L }�
��i8q)	�x�8����r�?���u��L½�Af%(�e�󜈔��q8���WU{�ߡ�?֤����b���ؖ�����Ta緘�lޣ�"�9��镦�M��u���D����}8�x�~����w;y�q�`J�!������:ꎱ}�oD�ln �E�j�M�v�_�V�x}a2Q�7
l��U7�t�]@�d�{sF`n׌)�5�������Ç-xqo��P$0����L��=�4> �|UE#.��-��[�y�oi����l�K�޸0�>���L����w�!�_萹��lOv��-t�uBn�Nr]6t��fYS��0c�Le��Ȕ�y�mt���4bnz��1zy������\ɵ��z�E1L��ol�ܝ8H�
���ڤ�N����gŧ���a��G��x1��ξ�����|ͺic�ٳ�6��"����s���A���nT�JT ��"K,]�S�6p��q\&5�O��a��W�k��{��Z
b�J� �&.��ʔO�U��f&��Kڿ2��;Ȋ1"�׵Q$N��ń����kf����G�*87�$]QY�~������Zn(^�uX������"�틨���Dk�����~����N�G��Q�����]�C�~����O��>#�B��Ӈ*ucS����)ǩj��%/�U7��j-�W_���I��x���I�yD�QӘ�x�tݻv�.���o�"�tX�I(è�F�iV�٢�0���NL���	N��8[�/+����~ 6d�G�P��)QS�FY�Kى=�����e��6X`��aQ+'p�{� ��y��ًA�SX���-R�s-�	�#���k�z�VUF���)zU�������ZxQg�+�
�D��\�E"]��iC`���(FΉz;~�{y���uP���2�6�����>.�!)i�� Vv�
Eo�[J#R����Y�������!kҫB.r.�d��vl<T��3$'C��W���,aE���Ӧ+�@����DG����c�c{���������V�@U���D"�{�u5Ek��*���pl$7���h��U�$�Q�8qɢA���S��6�;
x�� �.7Q>�);�L�&�4��0��u�/���ae��T����&�#��St[�}���<�v}�ݞ� ��J���xs��1+�Qs4# ֣}&V�w��Z�Vo`�Na��XU���!/��A�,5D4���o*�j_'��/�&�3�Н�5��
×1F�܈m2�����C|2}�F�%;y������Q>�"�<fV���h���m�mm�4���^�
���Ϧ������F[���s�&u����[ĞJ���7�5.|�Ws%F�R\��1�]��~��]�*{S&�IP�<�kPC�_�G f+�A����L�{�I�k7����
�c��xCY�e����h^4����I-���4(:��%}чTq��,�������j7��@��,�o���LQ�io�U �Pg~�Z��!���u^V?�t�>t��l�f�`IM�
����&�,MUh���4��qd0��^���$�Ԯ�;3��PV7�a�F�4���АZ34����(��J�n���w��:HQ��ٔo��#���V]ꪣ��cc���?�+_H�I�{�H*�r��n�(��(�x�>O6q��|���Ap��'hEYY9��w�|9^;�,q����'�#J�� ߝ%��K��-��^�Q{��r�Σ�^`L	a���#U[E��0`)�F�J|�}_kV�(��*����v����M;/O�&�����!}�	+��|�i0�8�Љ(3䉠��2=y=��b���o��=8+;I��\�;�(O��aj����5�z�P�I�i����^?��c:J�����I��xc�4yJ) ��:2�t�s6[�5�)!��x{�zؘhނC�\c[�zo��n놭�y���i����@H}7�WT\�nW3ۤ�V�Źp���O�J�1[�s�^��]s����k�-�>� P2�Q�	���()�h�]��G�75�S.O���>W�����	�H�`FH�({�o����Av$)�20d�v9�;�#�s���~�s�B�̌F�B���V�?.�}*��g�R�Vy�u|c3�q���tH|���f��u����`���mTL����`_��Ӭ�C/N��N��(A'���N)Ӑ�f��,|τl����ڷE*�Xj���C)�4�q�=�-H��X"�&�9���x9aa֟o%�=�V���?�D��uE�:Ep*s����!�}�?V�Oep1CC���q��t/VR�
���U�L0�����3��)#�����9�|)��������|�?t�<��=�$b��'�1嬽%��3�����������m��8T��o���QJ@1��@bBB��%�IJ�=Fń����衱@l���Jgm��ӥ25ܹ�c�Gaq �D�h|dqc��_�]O
?�|�|�t/��ZYj���x!K���po���*����$s�
9�:��!}���|����1����;:Z���c��^��4܆�X�j��G��-�վ0�����{����ll��ُ�	gj0����M~�hv��Ă;�]Oݼ�o���� �D<D���4��ԫە��� 5�9���m��{��B�h�`�]��˼Z�=,x��p=W�,�����c�V
�;��ź��c��������/D�Z���.D-*��.x!O���m�"*�0s�h����A��z�(G�
� @�;n1����'�ď}trhW����1��6E:)�D�5�)��Pk�j�p���BF�d�IK9U�r{{HX���S � W�-�&��c;!�z.�l�&R�����y)
�{~C�YPK�Q������W�+�Y2�jp�q�'/����l�Wi�����-]l/tA}����<�)�OC<�ߞ��
���&.7��v\�A@Ύ�L���p�r��k2B[���[�b��\��;U`�fl�����t��X;Iwm��`E�f�rf�Q�?����;�����H&�����}��G8�(��4k�/#���H]�ei�E")Z4��^,��̋K"����$��f�ni�I{���.A��c�GV�U��}M��=#�DǮ�L�wQ��7������룆�4Q�V6�~e���.������+�>'hX�ӿ�K}-��T�be�<�#S2�����P�1C_���l���Ȫ���@Vg׼)�z�0��4�M������qT7�rH�T*�������T�)��t�}
�͇9���c+�d\Ǐԏ�[�+B$n�a��Ui��r�F^��w ����Kt��n��a�T�Q�q{
�i:{���ڌ�t�8��S�~����URj�ll�9<Îqe���|x���g�H�a\��<��nm����چ�,���P���&!��(���Ԅ�	�Kh�� ���^���z�=/3�S�ӆ���������Y^Ntg�i���%.�u��-�f܋���n{��F���V
'T+|�<���AV.��c���`�fQ[��ި�2(����0�~Ru	�)�?�=^N=X�FuȘ����g^C������8}@��?O���C�-�w?�x�h�}���ߴӫ��|��Y�t5�n�T��3��^م6�����a�U..$U���)��)I�F6��2`��c�d�!T��-��t!-�A�?
Z�b甆��m��ۘ�C���Ϡ@�&����w�J��C�@7��^ŵ��M���hg�<IDO�������YF2~��$��ŗt-��)/3�ɨ��+�= ���n���p������*���w
	g]��B̷p��Z�P�|jLom��	�r�"� �?����gC�~e�)��F:=�[��*�@��uW���=^�R�B������L߳���~�(�-�����K�y�`0ב� r".�UK�X5�%�%B}Ih
�s����b{�b�[�@�A��,V�>O��pA]~\�1�.~��;��������2x}�֑|GX�&Tb�?��Pْ�@͔�h�f��&+X����.�����S��F$"�Ud��1�I��ߙ�>�J7�@�f�@�6��{�Rp2��������uCi�Ȉ���P�# ���&�������t���52=U�r|ВB#�I2����B�'R��������0N2���Y�����7�h+V�^KرJ����۷^�
���P�A�5�����m��Tz�~���
�3��n��}�9���h@fq��$OK9���.msL
��V�ДOT�?a�"�}c��Q��G?���KtO�j
�{/#Z���΀��{���o4jg�k��$1�2�K�{���ͧ֙p͎��{[�^��:�x0���4蠰CD]�}h���:�$V
=����0�$42J+���Ί０�#�tϻjw�r��1���$
F
h���i�G=A�D�fœ����WZ�SbF~$�0[8��2m��ޱ)�QL���J�n�[�� �0��^�!c۩'���NV��=sџ��R��A��u�|�~pG?2�.�R�M%�)��Î8�w��#v>�>*����`ٶƮ�W��+j�#k#O]5ԍ=��k���%�_��96Þ��YH�W7��I�~��U-�p�-=�̋9���ő���������5����U�=6�;P@�B�����ꈼ��65�Eh*C�N���F����	�C9����}Z�Օn�9|HQY�ӥ	+g�Q�׋���Z�]h�����W�&�B>�w����;�U�0���-�ʖ�)��n)���,:|���2]�9�|��a��7+x����e����� �6sK�Ӿ=1`@G;m&G�N2Ƭ�>�"b�qT|�)Y%z�ڬ���!��%�|��?+�٧��X7��� )���\4q�mN�&U�&tS���a:t�;�\MU�y$~��щ�)�#�H�n9$�iRuDއ �u�#��:�|r���)!��攤	 ��q�}��x]�`ڎrn�U1Lq�DU[�u �ˆG]���� �<Q�=�p.�)=���$X�/���7�y�n�?�� ���ߣ(�ɂ!;����>�5P���a4�?B���?����#�}a��G��(b���zFT�ŪE<�
,cڻ�1�Z��<* ���$�-P ��hQ��}J����~=��US��� �9��s��ڮ����]o	�f�5Dh�Bѿ��p�Y����
ć�m~����>�.59ʠ�z���~�DQ��s�X�����X�c57���L�V���|�a��x��g�C2��]�[O�o}����dFO��G:�2�ݶL����I��~��so��+�6�ܬ?��]3�p�r+߫���� �է��ʥa���� 2跾�\&��Q�˓�m����V��l��zg��Im��O�:�Ԁ��{[�����q��nRwTi��P�B�l�f��V����w� tR�#Gꋒ���N&��},��d~��@n���$�=�����w3� �GojD������+C���N7��'����P��z\yz�Vd��X���~��!#n&U�������^/_5n�'��=�\�(�@uoM�e�E�;�=�L���;23�3D��l6��QT@o�/�I ��cbD�UOJn�d��Z�
� ��Q���'>M�a3%v��'����BL!���e=g�{��Ȓ(v$�RJ��R<K���L����3Q]���?
\�F����/�?�_l�L���C���=|�֣���ϵ���:JPo���]�d��(���G�s�����޼,i�e�Ł4�uL��$X�f�ҡ��#�m-�w	v�x��a77�HSO5'����^-.�n䖷$���G.-Dz��-�H=K��6�	%n׋�����h�eJ,�2�F��Ř����%\���;k�8�f�,/�Ȗ���LH��zZk��T�C�F�G��E��C�l����	�!$���0����ְ�8~=ew�ǵ��<��+ y�iMA�'�:r"^Q������i��g�?�6�b��t��\�2_ E��7V���~[�v�T���J�s'���ᗘ6G�e��<���9;�%l���%M5��6 ��L����H��=�H�	H�+oi3�/��&��!j�𿿑���Q��yy͛TWM�n�d�ct�B��sʴ�"|������ɱ���i���xL��+ݵ��B��)9�_����r��l��Ǖ���%��wSs1��>ȩ��+����d� BT	����y۝n��D�O~�$����̒E��o�M?�;v�'��Z$�8q�E��?���z������B��OR�}i3�#�W�T�����8�8l��Ȧ��X��qG�RܦtC�/���S4��a*�Ȋm�P���g��"��ÐJل(hTwbr�腄y������b��8��&�ѡ�B�?h��
	P!X
�~Mr)�]R$e��Jd���>i6e��g�@���fՑ<��ؘ��=���qaW�&nԈs�7k�4�i-����-�JR.�����f�zH�匠���\Hח:�	���l��.��[��03ko��c��;��+U���D�%�LI��ĭž�V�"�T`���R�זǍ��m�8�6��(����яC��@�����0`�z�͒z%ޖ(q2���TTb*�2~L��pZ1ij���`/��y�����������_R�,q���)C�̒I��nz����5�|�/�{X<D3�,>7�Q��;���V�W��Kɤ�-��u�_3U�f r�����	J[hqs/,��� �)k4��]��9�m�3�e��M�͸ �eE��i;}�w��J�bIiY�S�7W��ЏM�����?�F�_sa/}�F�њ੮����*�|�o����y-��	O
��c�<��dw���ޣ��o�2��/Kћ>�����$a������|��}u(/�9�`J�6��f�?(����������n7�D�|��1�!q�����~���I�*��&v�= <x2O�LA! ���&:q��]ָ�&�(L�Sx�c2d�e��ϩ�3�S��'�N~f[;������z�j��o�6TW���t�������?T�Ҙ�ad�<x"�g�S�V�>&ڸ�Xa��"Y4i�����`�)�~���J�v�-8H/ї7)#%]2�����a��eK3�Eb��%���x�K޾��M+�����2Y��WQ��'<S~s���Z�����(�=PwgTV�T��M�Tr^��@a��~��VŤRf���!%A��S�7����܌2��V-k�v+KR�Ȋ��3x���O�{1|�U7�m1K�U����~�`��"-H\��,�!Oq���z8Q�5�)���<Acg&��j	}��!L��fQj!׉�#������yr}/���a��x�w�t����Q���*O6KW�Қh1RX�V��
֋NI=�m	嚞qG�(�ԫ)�U����ֿg�͵ͩ'EW�&�-�GG�N#�y��1�;�'�|�6����V�-����=���6.��6kz�t}=�ק/����4W�!�I�弄J���h���=���w�u'A\�<�-�6:2[Fw���a�iVA��Z��޺�$�W��?N/ �H(�'��g?�����5���Ů���蟂�?�s��q��qqD����=���Όj�sM3%�S( �o���?�u�=Ȟq�'S�§څ6�B����ې���2r��(ɵ˵��;LP������`��/�Ҋ%����z{���]�xX��W�C��&hw��W�[�-�\Z�f�	CW��#)l�J�I�T�D�B�f�Y9x��~C�:3{f���)��$���$�ꀆ*e���Ź�%���\He��Z1F|W������؉��x��r5�%��p���^�^����{Ĉ�9T	��},�����EB�Ԇ0���#
'�PW��p��(��Ep {�f��(�A���JVټO5��ߑ���� B�{x��G}T�ᶃܲA����!G�B{��@���A�.9���d,4g����,_�&:��ճ�j��gN���m��v���	TQ��-�j�1�غV���x����T�Q{���;�n��}��:\02u/��-,(�����lw�8��P~5�D-e���,�E��#�F�v "ݗt�r�N���H})X�H�P�껋�]N�R���3Q�?��-���c��٬+��>�
Ժ�2���'4z��|?H'b���+�珠]��@�$^��3��W���T�c�f�[|"鶠C�
j-(�q�7�L���c+���T>��byͻ��p�V��4^����l~��s��(�P��spi���y����|��v���K��IG$=�@t>�P^���E��@O5�_�Tc���˵e8��^R�̷΍%�m
y2��#=E�n��X9%���IZ�G)}:�ё�(K�ӭ�8*7S��Z�|Q(3�B?����G�t&���kj�L�,�]}9^g�WSN�����b]�)³\���LD���Nu!���
�"x<���/8�G�R�lf���]/�s?�-��p��O�Ӝ��)OL���[���7C$-N�����zaΕ���ƮG���Qk�:1���Ѣ	��Z���)��C�Gl�Qx��Z��b=f��ٸ��r@TȚ��4���+U�NB�H��lc����	�Q�a���:�� �BYQ�K%��WW����CZ�X.
N�-Ң[I�_�Cr+��]�	�+"��}�A�9�I*�8�ޏ}����и�]	�˃�pS�!�M��l��[�� 7�G����`�JL��'�桗��7;6�o��O,�'s�[��˭_�N�[���Gǂ�ul; D�! �b�;���e8�^�,J���1�[��h��p��M����<�����T@�J?a��EE���Љ�ʥ���Pl���u-J��B�lC �qd�>c�� ��Q`��H�X,�@���J�]��>p�0� �	�bu&4�N ]t�ǒ�h���W8�6�]/����&T�Ԁ\NP%�B��������S�)�ux�qG[��wGH�e���I���v���h��vb3�&|1�l���E�ih6�KY�Ȩ�����R���s��'�X���T倆���B���D �+��C�����;���Ϳ�R`�WM	"���^0�Ő"Dv�;`-��M���#hv\|��,�m8}��0��Ocg�b���W+C _����7�Ƣ�k�L�|�NT�W�
��}�D$7W�uw���mb�6p�H@��k��������m?p������PϠ��pB������ �Bc�3���7h��.�у�+-���"]���T>[q����X/¡�VFXOx�
����?ʡ(����O��1��le��Tc"�p�8jIM�t)���E�Vq�oQT�5N���xm�ƗVBql;țV+߬D󉢃��w{,K�%���ꌊ0�]]�V���E�55�`T�f�p�4�� ��}	�QЈ�)��ʳy/���IyC�Q1+>�>���Ź �"������uNXɸ}΅KF�NhA��,�A��� �����HrG�vw���A,&?�B2G��o@G޳6b��^�f�4��׍Du�5��/����hBƾӎ�f��]6�c8t�_;��'|�Ȯy(
[���7��%�`j�i�������BXd��T��#O\-�}��b��9_Q�(5/E�wq�&0���z5my*�o��DzZ�m6�>R�����8�jA���|JӠO�ɯ��\U��	��#6���2�[��T�(��@辎�t�ryIv,&�}��ܛWy��U*|@`E���g9��єc�OG�-��}�x�e�q(���S��\���%��9�=��wɔ��iI��Nz�pOku��Y��"���D��_�u�?��t��ѯ�rZ�sU]R!O�eC�IՀ�8ep�'���$[�䣵���3P�8j�9DkǇ><��X��[��'�=@�S�Id�ެp�m�7����]2����Lt7�Hk�o~b������
Y�4�=�nL	�<m#n���}���d�+��3�@��1JX���x�����5��Y�QQS?�ke�����t�V_�ij=Rc�-����C�����*Me�Ywb}��lC>��iMM�WK�
!Y��IX0�i�B�0�o^O�[�k$� �Q�)�	[�8t���7�
�Q�TKJ�����/]��a%:��G����
�4$�޽wlkR��I2A	A�0�5�A�s����?����k�\�Z�uYE���#�Ǵ�so�X[����p���g�	������k���e]�5V���i�
xd{E���gW��H5"��c�Y�
s���M�'�;��6Bx�\����Ww}�����M�1l%mR�@80-,�Hħ�?�b�a�����M�|��/��nh�+mB�_ep]�'m��Y}��g:�� e0�i���mR�![����h���9��\�kFZ�
K<\�I�m��~��'L�:��(��zOч?��vz�j��=�[�`�䔍�u�9����,6꼃�b���4~Upd��V�'��h��ۭA����!�'��2~�怩�Һ�ƩDGUM���-����5-8����C��Cl͒,��i����t$��ƶS�t���̸������nYe�<m�O����5����"=9P[\�<���*��;��5-���.#���_
��/�����E���P�h!�2��#<�`�z͌�Gp��q�a~;�Ol��P����7(�spT����𑂐^��XL�*S˕u�!�)|^��}��w�_��k���vK�<,���Vg�Ժ�����^F�3�ug�z4�.K�@�Ȝ����G0��|�K(�
cOI<�Q�2��YV�8w�9�5� )q3n��
ZZ�	� �Ja f�������x!*c�F{�*ǃn�]g�BBW赋�}V�h � �x��}(�,8R�<�X���]�?+&8["�e
�5="�Ѣ���s�"f�X�_A���._=�ޓP�FΩ��δ�qsb�1YISk��S~�����6E������߯����������E�q�X��2��|S嫩��������)̩:��%��i�K2�n7��Ϩ��
$�L��׼�|C�_Y
���s���W����3�h#��" ��{��8�^��[��:^��N�2��#B�)cحĊG�ַH�u6	2���h����b��Zr� �c�����G*�a.̷�}�L�����M�Q-n�r�۪�xÜ4C��p̝�H��#��l�e1&�|�I$��;�5�R�+�a���@N*����w�(�(��=�]�y�ʍ�p�I��� S����w���4��."'�,V�(�	S4�q�/Q@�B(����a{���h(�u�f)��Z���f��[T��$�}֕u�8;^���y�6A�%c�7�*>1g�c���mQ��WeMh����PJ��V͠�a��7��<4Ow���[p�͇����'�NeM���{T&�]�c��,�;��/'~�!�hz�_e�u�
��+D�b*��\ dj�l���[� �#惜'���'���L�5�/�a�OD�l��������lQ��m�GT:�	���x�Ԥ��j8�p،9��M�kwd�~y{����ƍ�®x=���^��ũ�U�+���<V�b��"�=�,�y���������7�9���[�p`5��š-����"d�3[��f���6J� Ѻ�
q�8��?��K������T%���˯��M�&�H��d�%����N�W������΁�;U�l�I��2ǭ;�>�j�`���Hz�s-e�{p� �U������j�r>$4
fJDσ���c�s`Q�|6E�s��Cg���a�@��B�$�r��?�
����x_�l	�B�͉�h%1���GH�iwǩ�C]�QUw(����I��-��9�E"���/���U�oK���`�rt�H�y-�d���y߮�<�n��5�sW$���Z)#�!g�hvN&�����QB���ˇ$�"����x�so>�__+ٺ&��X����ۻ�^~�B:\*1��G��N��*4-��2�X����e;�l�,��f�a��EI��7���MUuI��+��_ �;�j�_����gW��@�pkgo��1Zo�ӎ2��V )kT_3�@�����\�3�T@[e����j�kݪt-T]������cVvl-qm��7�P�˖�횪����ȑn��<%��o	��)5R��A�ٸ��C��, 4�.�&۷�%oI�	��~`�7jG)U����k4U���2ٳi �P��	�ԇ�M�=��H�on$�`v�ݠ!4� {hG��̏a� ����|F�ZȅJ�⠳��� ��}��G��=M��*U&��[�Օ1J{ʂg�+�G=���z�L�4�b����G�ɐJz��	|�g�;���x�e�P����'�@g�ltQ� �>e�=���I�Ԟ+ԚvA���Q��!o�g�ڡ�z�{|2ţ����Zջu�u��5�x1��I{8a`���x�I�NA��.��k,$bbdj�rG	I�} �x��P��<%�ז�;Б�>�O{!�DT��k��* VBs�R�A�+թ��pj �������x��S��,*,&a2ȭZ�����xGJ��8ۥ~�i!�
�;�)׳��[P"V����S]�����7�0Sء�To���@t{�����&���o�`E��\����������&AL˖P n�ݳ�FϷ�ݨvU��?�w���:`C:�]D�x#��}��v��*m=�����K������a�=��� ��݂�q�߭˳q�%��(�!�:_vc�sx=��ؙ����8�		�x�R2�$,4�_�ޱ�ł<Yy7�IS�	5��L;;r�-��PG;���*f;<.2.���`]M�P���=��@8,_6�^��񂠽�d�8�~�������iI��9�I��jB�R�phh��i���lj�(}08lH��>�Zp�h��6�ʁ�Kåp���)[�]��]��	Y�<�;6h���K�<Ȝ�����j7N��>7P�:L$���n� rS����j��i,ԋݨ���J-�������8bv���7�����?�����f�ԕ�N������YT87�������U\�aؿ��f�˄�{Si�av�D(��@�����!�&�۩��9�팜1n6���67�pS���N���h��a���2>#�ng/����_��h�!�y���\n�`�w���Y���
;�5o���h�$1vX8<���ԯ(L�U�"FS|Gf��������r�����v��1��_��\�Ծ����?���k��:3�Go�M	�Ly��d��Ηrw}`� �c���� ��\�{b74��V���٩D������G�-��D?�i�%�vd4�-�nh��d+��ǌG$fK�6��.��:��)o%��*��`�ԑ6����k�X�u��g�{�'X��R��a��rH�5�+7w�W��(h��T�S��2��ɛ%4-����x�J����1-!a�������خ���#<T��Rp�1R0�`:ә�Z����,-�������ӤQ����Nas���D�Co���M$ƼA���{A��
JΧ;&-H����Q�#0����R1�Z����T�6v� tԊ~�m8�y*BvE٫d�N�v`|j�NI
nf'�����sY�z�����<�4�"�1;.#09:j�ʕ�Z����T]�Pψ�z���	�������s�V<�Tp.���E�~S�	xD�#.�,���+�q�*+�qh��G}C���[�r�>R�U�9}�Kh��鄲f�ܽ�R�nS����l?'��9e7�,���y#��#VS�f��JZ���_׽ک�$������5�����g1�;c�57��q��qY1�2zޝgL�����j ��3�����{�ί�Z8�A�o�H�B�V�YfZ����F�-a�"�V2�⍒x���&�}w���0C���5��PT���1���sp���dN��w^^z�v\��~J��K_U}��Hm�&�!9 ��>F#[���A��9��fM�:���q�ЬE�X�Gh�H	��"�=�К��X:d��)͎�M�y2�����*�HV��gyy����n���GX�sÈ!+<&�&Rb|]�DNh��f�~�C�b�hQ����=&����P93�#o����h�1�_�k*�6,fV"��}B�N��jo�ϱ{g8�#4��eR
���Q��׀�:Ku^��p������ E�u��3�����S��]�9�>�*S�!�+���w�
��30&�ӽ=Րw�����c�\��
CCr��lh*0cl+o�]��3>E�i+��o�4n�ZWt�E�6Z�R[2
���p��R�+d(����Ǽ�WTe�B��EO�?�l�����A�q'�fae;dc�c݀����ʄ�K�#U<?/(��M��5�!����+;T�S��6�-�Ε6�����{5� �~�:�@���2���7�V^�>�X�wiə]����KSj3�I5�*u,�v{���a��g�����|y��2�G�?�(��)����֒��U5c�8�I�<ل��a�*k��=~����0�d���{�X<���e_�ATVb:����.����
�a3MM�7yQ��}����K�=j���C�6#�ɝ�j������������*�@�c/y0�J3���8����u�DyO0�蔏<�0IqT�⩸a���P���#E��[ؔJ{8��P}��߬$�"%Vh�&XF��}3b_<pcE��aQ>H�ᕽ��$wn� �-eL�$���࿬@G<�;+�r���R'%ͅ����(2���6�FQ,��g�v|�Ї/3�_�w�Bhzo*��t�Y~.󗞯$��י�����0��el�W	�)���u��j�'�ǹ��a��3�Cݮ��X�K�:��9n6 �Q��(��,g �"�G�][�d���ݮ���t��!��Pi�r'��G�V^Å>�E%���$	����~���D��O���ɒnT���,�ݓ)� 	b�����~��������ܢW�w觷gDv��	ϤP�?�W���'ꎡ)g(:�@{�BU��P�~T�tgo���wZ/r$��R�C�w�����2��7�Utf4��v/E<�0��]D�Jx*٣m֭ �n����ߏ���TGD��U��̈�����F����Z��h��w��Y\�ܟ4�@��Kb瞅��)E*����r@ޗBO��� ��4�o�>ǎJ��'�h��V�C�K�m^K:qW	�bK�:����R��
����G"N4[�H���2����A~����v.�`��uT(��[��~������EqV8��H~˲�M�&F�f��X��Q̈́R s6��k����Y8�>
tCL����,�Uٌ��QeD����ø%��S����T	` C >��h�c�1Hsp�����d��za]RTsŵJJ7L�a�Q`p��h����0�{��A��n�>�~?���O��ڈ��@���R|�����쒄�B�I^�=O~X�	���1 G��ӯ�sįB3�e&���l�q��E��ՙÃom������(���Џ�N����!�a� ޵�U��7u�����|"�fu-z^0�xF���)G�u1KS*������6Y@��O�v*9���YC]�"�^r(6�������^�������A��~_���e���'o��P�#�ͫ����jhэw5󰊵L*�����	�фv��Ұ\0m����X@c���=�}a970FRj
�ĵ �<�����_���y���N��jO�3{����nѵ���?�`��P� �w/��:@���j�����?B�����%a���ϊT3"�
P��ap�3�8�Įb�����2B��R �85��\Z�ܶy6w� 5�8�m`$-6���
���(.4����yDp����c�VJY���$}�"�^K�B�-W�)�d���]p��3,�]ƛCJ���[�Ǜ��kr�����~��D�*��ȏa�g3��Dk�V�m��؜AWQ_ŔY(���Ԫ?����^��֌L=� 5�5q޳T�c&,�n�Ɓ����x�0I��xT����W������vu`��a�9���a.!h1�:͠�	c||����V���]Q�8/A���N�o�ǈx��e&UZ1R@0j9��,�`�=�F��X
t����/6�\!��/�>ry�$`��A��$�W>��޿#%�K�� D&
8���PO�'���;��Z��7�~��6� ���4�t��P��:i-pp�~����J�f�O���hO	p�.�ţ9$�X���' �w�pDs�� ���9�2��&�=sۭ �M}�;����r��D���Jd��qv�B�f���3�,�������`���L�T��I=8μ�Uw��D��,g9��m��P�����s��P*S����D
Kͫ"q�@������e�{�<9
v^?Z�`�-��V�P-�u�����k�����'��v
� 7�����1��`��T�?�70�i������������4��Q���(r���-sC���`���gk�5�lzYD�B���i	���չrM}1��Ď�6��W
����.�7��ϰ�)�*���/���PE��?��K�=:Wd�pݱZ�����\�f��5�[E)�C���S�W-!���5���hN^dE��*��&�/��F�@߁VC7g���xc���}�%���"�ե��P���`����Ή;?$���/��ހ�h��#X� :DB.�d�l�c��s1ڛg��8����ڦ�ZM�9�4�'vQ���!��SܖH�h�ᄫ��U�  �N'M�^�r�R)�]����F��������T�A�q��w�N�S|�FSM�[o{/;��p�cK�W����Z`�G�t�+օ%l཈���9��4z�A^�*|P�D��c,SFյ<�R�@�������r7)���b�j̔�{t#]�N�pO�ؽX	P<��a��i��as�k�M�f�,�<�r=��zX�~fM�l��E;b6�C��rݾ�J^N{����^���UO�a�~{?�ß�s��+C�fe���^�����UM������H�Oប�Ǣ��^��i[�pƿ���� G�	q���2�ql��u��͂�4l��N�̀�S����tϟ��è��q�4nr�����<��.WM�a��z�kNe�E���G"Z"[�tݘ��]�Q��yBU-/ݘ�B؈���0���������?4�Sڡ�De��;
�Y~3Ҏm=�Ĉ�֘�;�g�����q�5�ͯ���r �)ԯV26dË�Kk��I6��mc����\k�ӆ;G�7 ���E����2R��lFaY���!0���ֆ�`��]��:*�m��T�f	���	퐿�8��1�}=�ע�A��i�*'����R��G��ք���������yu4�6��ǆ�gu��!D$/��v����eP�xn�E͇#�1	V��(�v��z�DO��E&�e����4�d]<@p)\B=of들��s
��m��ћ'�7��p���fM�$��cd����\z�6�n���j���6J~^�uRƭ��m�Yu���k�3�cr��lR	Y���R\�a��~��f�D�p?i��i��eZ5 (���|��G+RBc�����*�B,@�Z�2�Y*ֺ�=��������ځ����_�p{�аMNd
C��@*LP3��W#�Ԥ��VwS?��X��b!�q�6��X)� GOҜ(����59��Q�a.]ݧc ��:��C����.'ʣw��[h���o���ORN�.O5�B����uKz�V-6Qy�� 7�0o�X�ɀ��!t���y���qE`5C���>�[��7Z�F�.�C9m	�c!L{:Z	+/v�W��5��3��Uߓ���Aa��@cNJ/��{ܬ�S����n�\5��ס�����y́8yM�Hk2c����M�$tt�l,�������{MRD��GtG�&�7�,$f���v���jWv߅֔7"�k�
�;#�P%���W��z��9����{46��c@��&fe5�1s�7�P���l8��)�|��kW ��^W��h�a5�Ӈ�� 
+]�/ש~�b���.�g���D�;u#���қ�㪖����S
��(D��IWf�H�B�ǉ���<�-.z�b�Ђ�OO�b���m��0֫c7O^�xҭj���}���c-��X:[w�\ݍs�8֛��aZ��gGˤ{v��f�t��;�	�Ɋ��y�����E�Ƥ��p����h�"
zC�k��T�[``_�ق5���L��M�Z`k�s���d�ߓ�U�?Ro��<��~�n��*�#�{!M��u)$����I�u�LVe��fa�
I;�JqUb�c��s_3��n`����%�&\��"�L�����|�����D:�.r?kǗ�@%��k0ߥl}P��9M�G�俥G^�T��rK�@R��tb�?�iB��"��1,k&ڲ^�z|F�����c�R��\\���@I�K��}��h�#wG�)��n��b�E=v'6*�tL���˯�¨Zָ��M��jһ7'�E~zwL����)y�᫖K�iK�dK��L���ް�8j-G�}%?���j���O*�͆�&&Xs�P����+�����n��GR���Y�o�a���e8��_�
�;�(RX}�����9�,�|��s�/!�#Fc�"�����E�bG�t��]�RtT��vaC6�����.�8Wg�n��j�lh�a���B5�D�
ǟ��|��He���EkX�q�J���%-.n�jn�(����A�d���/<���G���LR�b�I���x�]e�&�����a$�6'���6���tN;!R������-!|�6�F�^����d��4���z]ιW8]�?��1�w�p�[Vynl3m.*��T��Ѭ�L�Хw`j�U5iF�BY�O _;���7ˢ/��%!�ƿ��2ِtTo7휸����\l�������r�8�(�v=��@J�Hb2��b4�H��r�;&�@-�Ԣ7<�o�Ö�x�����2�bJE�<�%����ݒ��޹%"ʋ*6�"N\���F����]��a�umG�g���8r�Q�}������F��n�4�
 �֤�KPTR�Z�d�7�/\�B������Mه%��[@-~k�p
MR�t�s��;�Xwb	���##4��3�
_8Y
�;�ʑWPUF(�O�L�b6&(ؘ#��'D�ɩ2԰O,!
��!!�մ}��G�j�h�bR"]��z�ү��E�@���27_g��[����P�}�D����Y�Uw�=A9b�����-��4�M`�be��_����]�*g��jy�%���&7.Ҥ�������QC��j�4�Y����[�e9ՁR�#��0�Ϙpc�m��`O�S��u�&��x*[B��\��o]���e�K�7N7=}D���#�<8�(�i�*�3/F��5�Y���ׯ��1/:h�����$�����D����v�����h�`�C�2o���\�^�<�@3��V���G�i_�R��%DvTqr�eݺ�!��5�����u+�ӦK_�H����@���m]R7�[�[�>����.�%�J\N�S�� �H�(c�K�醙��!�J\�9
�����=e㤦`|,-Þw[<��M܇�eA��C���SŅ�B\�����	��ȎA�����TM/�4�6�y�:sg�*~��ð��r��8�EZk^F0,>��z��\�atN�9/y�D�Q�|���ק��Q�<A*�b�	�����F��m�Bu'*:���(�=���o֯;�f�Iz�1Yo�H�1���˨/R�Q�<Ǭ�@����@�ݏ�1u?y7Z/G�٦qm�	�v���=-=���>C�g���ܨk�ۑ��2#8���Ch���s�8�2��b��#b�r=!rK-O13p=�צ�����}����>N*�It���,�5�xA�,Ț�G.x2Ƅ`����(t'�k��2������^j[�h
K�xrk&W%.l2��57Hb��NP3 ��t�������Q���-�&��.U~�IVװ9, �O��"��Q�4�/'v�۳펷�g���L-��n,������u~uYש��3>Bc�x�W���_&s�@�V�--s�,5�lt����>�ӈ�#|5nTݲ�y5p�
ܳ�*�[�0.H�2�Й�m�sF��:�t^I���HW�wR[��y��'�-[��$V��Q�����l���d6^�=O׆�
%�kX�K(Ӻ��c��Qv$K	�r���(=T�ƣ����mM�?9�~�	;V]�5PD�A���m�=�7a��C��t�u�|�>I�
ӑv�`���1GA=P�#����Gcv�q����w���<
����.���Os�gb�cF!dR�H�U�E
���	_���� ���92g�_��q������[Yw9�Y�"2~��z���]�F=��DU���7!�b#^�8���	�W�+xur�>$��Ş3%�B-�(\�j�8���S����Ka��dR��L���WCs=����>�#3��e�L�MN����h|���$-h��('�|K'������͈4ɏb�c�`�oV �܀˝$|��٠^F,���s��}5r$Vn<q�t��YLt�S~4ę�X|��@�m$�"J��u �:*��� ��v����m�Ǜ%������/�&�ܺ����b�䨣�I�7T�7�y�@)<�L�\+��Ld*�@��c�����p]U�"A��J��v~�h��;E쇿 ⍱�:��0��˨ى@{͞��ܘv�rae�{��s����E<4I��*���8f��N�� ]�[��6�"��|�K</X��ƫX�g�&Xb�Dg��qF����A�b��Ty�0���q�3���
m�ys-��_�{G���!D�o��#}oQ��z���n	_l����������z����<S��H�AQ+/E`	�����KY�â����(�}���!�y����?�����n7a�����]n7���(�J��Z��n9% A�%к����b� ��ܥ���U15�'�8�l���|����}����&����	�������Y�K�<�x�S���I��=%�b��YI���$�)qO?)>O�����n�T������aeH�gg蓴����\e#<`���t�8�µ�U��-R#(�Y���;Խ�q�S`��J�� �<[�6� �A� z�\�����U9E�XmT<m}��M=���וptm�=�xƖA�� ;��th���R�T�Fd�~��)S_S)�LtW���
�Ʊ��.Y���������<�g��Qw_�����R\QF� ���Y��Є�9��S�%�P �����v����`&��y[�0�+��d0;����&�j�ô7\D�xuM��a���������z5�XE,+ C�D9�7��� ;��p��f����´kP�u6Ly_��u��m��j�}��P�;�;>7i�N�ɡ�-�}ْ�m�D�m*Q,py�IjkI�x�~0�vt�����L~�SEu�ͅ���`Y��SL�s����|��2Z~�"��v���f�O̷���*�ӚK�����2�R�V���{y�dǤ>s��өy5�3��ǻg��S�e�wX��:���x~.W�wT�pR����o[�T���fHx� 4����0/���跬�:�@У�À�Ҋ�E�-��j�g#�jl��}�?z_eT\�Z1�����C��T�#�:�JM�Zq�Ժm���K^��;d`�-7���S�"@�'�KJ�r>����BE���%�&���~���9����1����-�@���!���߷���ՖV��;g�t��uC�PN�s��2��>�zy��67�"�l4�Kݝ]\�i�U4BUEa��Ԑ��)�@�c[%H�D��^_&���������i�.N���Z������v�qʃ��~C/��}ډ��}�e���d�b��[��4:�	�@ebD���>>��X1��f��$�C��c^������Mw���.C�Y�[-�����w�E���BL�?��m���E��h+�8�26Z�]����b��W���FC�Hl��R�c�%�A������6�eFU;���ζ�u=v�A�W� �7H|��� ݔ���X��|9km@�lcp�����
P�o�b{��r�����c\�n{�{�D�l�V���&�s�`�:#����\m�M[_�n�̫^��sQ�~E�*�⠂��͓�м�F\��A�E �_5��jt^��;�m/`�e�9�L��M�[�ܴ��P���G��9��(���>l��5��͛����=)Y7��3�FXWN�W(Nm��5�����F!��bV��Lν���HmSJ=.*�7�m-o�������ͼ��k0[���B|85O+!0�Q?�{?�P�Qge�;4�\`~O%�" /��8�v��<��}7%y��Rֿ�0hj&0�{�2�����8Q�.-Aq�kE��:N�HJ�F���W���,Cc�-�hbU��Z�D���U,f9ۄ�LYً��M�4�����P����т��N��U�JH����7q��%N���˧���wRo���H�Ojo���{��0�Z2_�*+���A(&{Hd^G� R`��g�̬>� ֚TC�q0�Ü5�ws
KV���^O4"�&^��"l72:F��,����ǌ,�<���n
@��R����y>�ZCeF©G!d"�X7��]�f�C���C�r�Y�5��}�//��ؠ*��O@a#K(�t�����lct��dL��+�L�y?e9��� ���:�x�Uo�=�dO���k�s{���\���~*�!���9��X-k'��!�q>^� �)�gj@6;6k80��?B.ۼ��7�.ur�B�-���S{9l����{�U�M�tg�`yQ;����|��L|��S��gy(�ȼ� �P�H�~�fUv薟�;׭I\�����҄�M�
�I\{ϴ�Fض���N��HҔA�~w�Y=g����o8��r�5WX�Ǯ<g�/�Bet��G��@d��_��%b 	��>�k�����#��[���@l�=j�QSjL��<�!E�.޻<��$��mE"�M� ��s/�)Hn1�Upt�u*�#<B����TR{�E�g� ����_eN�`��r7�Pָ9���\���$�U=t�_����:a��{�c��*0���ΩH�U�@U����4�f��)I��i!9���taUA�򷩅�B��' ����Ks_s�@�x6Y5+I�g�M�ߘ׶��O��#�UZmJri=����G~T�P@�q2�[��'�3��J.������������_[�h�P�f���M�\�	iǟ�+�Y;L�����f�B�Z�;7���W�^N$+�E����� �:�Z*���Ҝk~�d�Ò��dTѫ��>��o��e+��e��{� ;�gG-��KH�J-�Q�LLቢ��A�ʾ	2�4~�y�_���P�ʠ��>�ν[���d���N$/OѢ���g�OK0̳�,�a�Z��,bA��aŶ�`�2͉�>4>�1kĢʅ�K��}J��[|�ZQ�>����cG�:������)������&�<M�s��'ڶ��R�Ъ_Po�s�m���;�D�l2�6j!@eS��/����4�G�v^���Rq	:L�D�c^��1�[x�����{�l�>O���`���(x��q�&�F����k�W����P��/g��������ک�u+(x1t�N�F*�Q:�~J�������A������	��JtBm*��1������*Zvw�i�aa�)�D K��ǀ� A�׋�����W"Ǌt\R }z(w�%#��E����@-2�N.��*7([��&L�F?d]\F���5Pj�9a�[����z�����ש�.��Kc���$�U���E�3{R^49� �]�{�0�ا�D�M�l�3о��`�e�&�Ρ��7�d�q+e9A_;�`�h��r';oԺ�c('�k��V��|�]]l%��{ZÃ��^��U��O�h���٤�+N�,-[V��Fq1��'��.G�-�zB�|â	��cX�偙������1�z+���,��2�R���iPX���Q�4D/�%��Y�gZ����f�JX,	�v�)S�q)>�K�y�i�&_����^�{��(K	�>�Ub��Vt��죭�i ��jUr �5ol-�B^�o	n"�j9_Hmkf5���yT���RL��|�C��fS�wB���������Ћ�
o ��N4*��<n�z')*c�'^̴�&K��4�;�j~�3�e �8B+��&���v�^���x�|~�ߨ�'������$
�5Z�����B�Ʊ�xx�-ӆ�V}��q��E9@�t�G~冭���!��FB}�ٜrG��,_+u���nbaҜ�)ĸF���dƱ�1ٹ�����$�$�Uk����Mou���M�8y%����bAp,�!˄�dPv�2�Z�8���J���a�"t�-/f�����ի˙(�ɸb%^�i�-� �:�R���~
���Ha�nS�<Z��f�`b�7�Կ\�4#���@��g�K<E�$i��a�n+]��}�Wٳ�z��TA -���<��W�p�?�!�lV��x�ǈD��00[L�j��� s%lA2''خo-K;�hD��ŗ~�'���xhg)���1č�Z��f[�sH+�-Pt�il��V�M�&:՗��w�������}�-��f�YINf�c��A���9���^�Hm��	�$��~<���V����z�/�JW��rU
Eէ�����t��w������L����n��#�E󯤌=��
�$iF�y_�t2�;��$�K4{)�wS7�Ҝ��fPX>sZ(���#W�l�����A{�ƣU�ւ	k�2ciA��/n޴$R �J
<� n���j��$��):K���ݐ��o����:Uc�G�$T���`NQLۺh�7���m�Y�Qn!��O	=�QQ2��>��lav���O=o��Y@�P��	h���� �)yl��yBC��"�at�VH�hB�v��K��sY��o�@��?�Q�W��>dx�^�*�3\SW��B�+�Av�� �B�C��z�؅�|���=s�/v�Z����� ��p�-���R��N���5�����9ǟ��D���&��&aﬠ�)���顤 *�6�ؕL}�br�*r�N����*7&��GwG��lݛ�42:>�I�]6�4�,K߻R1!��iJY(E׊3�Q�Ⱦ�9�!�R���tB�t�$��B�$���N��VdU2
���	I�&0q�WI�H���5������v��E(�L�)��(� �o�w�wp�i���p��Sp�މٓ\j*���C����s����́6� (�W��jYM�oE�g�3n�&�)�NUe��3xo�.�Gk������Դ��,*��rm�ʗ)}Xhfݺν�e{�{���t��6Lhg-�%y��m8�:���}	����Q3 ^H`R����T��"7ܤfd����Pyjm�}$��2�B�G&��J�������t0c&N�I�\�S��a���N����aM��o{+��\5��^����H�׿3�/��2񯰥�5']���\}|a���ZCX�-�G�*%�;�S;�L~��;I����*�Z�i���j궤ˉ+A4��xN\ۋZ����mҐ�V2V[�C]��DF��B�E��L_�q�$*������'�fmj[�c�uGY���؁�&��X����=Ȉ�P���W��hO��@A��rCv@�GoCN�Ϙ�4�1�Ӈ��rͼz����v|��-j;� ����T(����o	.,ި!�1���ꏷt>�,���چ�:�A�`Zp�vI.X������ۅ��3<�[x�>ɨ\$cռ5\��3hpǗo�X�Ƶ9&�8c�a+�<U��W�8A6�p�h���Y>���i�Enz9Cí����a�,����y.�aD?��.{����r�R��F�����J\�ߧP�]Dc�.:0����ƭ�,ɴY�
�@=/�nGGm~���۟��Ug~`6����*� UJ���"E��B �m\�#2s+E@t�<6�K��3�'	۩�o�hKD�ڒ�+��/ �ͤ6I�y�����[�Ì��ϽiSEK��+XO�78���g�@�J��a	#���Jd��&\o؟���)�:�8�j��k��]C,�9�S��!�-59+@���HY�I�jAd�^�M�m(e���ص���5�Mͣ�?L�G�)gm%<i�h�f��a�b�Q�նc�YVg�X��!�(��o\��b� 0�B��z�?�)����HP���7}%.f^%2��Eny���TJ��E�f�Y�o�̀k�O���,m	L��+&�rU�(>`�=�G$�
,�o�� R������'��Xf �-r��K� ���� �pч��\���3m3|�D �����fȹ/�n`诸���ь`?o��%�7�O��~t�n��F�bTuG��.t.=!'�����~ا�$�@��2
���������ד��-v
����.�Ĩ[l͇x:�:����T�Đ�f�GA�fN��m�=30F�R��Ѡ2�����������n����|pؗ�=d��8v�0�^��/�ϭt��^j��O�䄴����V4���R�%S��
�R�66�#P�x,F��"<�v�W��X���5
S��ղ�/��X�*�UVZ/Ԓ�a�e�IrlA0_�Y�?+'�9=�㚙f�$_�����lM���5̼yr���F�=d
�}x�&<�>k��X�[MT���X�zq<���z޳n��`�,��!��p,.۽��L�^�$0��duCJ\�A��~ͺ����;�=Z��C�a=K.O���P8�(��-U9E�o4���th�2Iɑ��C�#�V��|���4�F��v{�ˋH�8U|]�G�l�a^yf�˘�O?��\͝�%�IK<>�gӢ`T����7V�\<� �J���Ȥ6�T��D�L`���+�&�{�C:��.J�s6w�?�偘i �gI����Z�'HJ�*�L&�B�Ⱦ x�랪�����_�4l�p��I���1׸����]���Ԩ��މSN S�x��Z�'�D�4���g�Ҭ.�OV�vx��sz����`5K��+-�� ��6���$�`��
酐�,*�V��r\?�;/�]�s#���� �pAV���|���%�c2ʓ���t���oa�s`��tj��ọyk�x���~p�q�>$��3��������c��`�=��S{N>�2.:K���QP8ݓ�-��#�]S�	=��e������, }H*�8.��٠4{K	wXf���-���`%sbVPb~���c%��R7,�Ikq)��!��u<Q�£��Aq�R�;�i�e�th9W���*J��>�S.*E��oi�.n�Ѱh{��F���$LvR%��������Z��u��E��b��Iy�&w���'
N<v�����>~v6�*	�f��0Uұ�{�bÔn�c�}#��jfN���v}���LN&L�9���װ�N:w�S�<ZM�[�{��,�|'{* U���N�3|�f�9�X�l?"E�&֙� f�'䝑���a��rkYH�`��*���m��
	��[
�#)q~����4XU��dJ� +f���g͏������� tc㜄E�A.�퓴�4�	5�@���>���I�ݳE�d|�g~��v�]u��h@�zK]�oؔ#N�#�{
ͤP��EV�{+E�\�%�z�7���$d$Y+OC`��/��wj[��IPZ�%�=oj���I}A�����ь�JA���~S���c��>#V�}���S�'É�D���«���<����ia|LH�{�I�5˿vR����"-�ڰ:W�9]s��=NSI6G�Z:�=�Lޱ�ƨ|s�E���a�e/���}�-2�����(��l��y�waR���� 9�B"\�x���F��-���!H���:��z��5�����ۉ=�Q�w�Fxn#�,9%*T���z�� �+��cF@��ɬg!�,���P�Ռ���{��[$ud�8|BL�F���R��������?�zhN����fVy�jRּ��|�J!��{��@@Sy��'�����i�Щ�br��,N~(<>�bA�zx��z�=Ǘ�*�k���fQ��x�Ue�&D�5d�=�XH>j�#>�V%2��1�aM�$��𠲂�"	�ok���j�5��%а��,��[�35�J���}0�X���Ʊ�L�b��Ҫg�U��ԡU��M�}�@�!H��U�7���<���2"P�cFQ�6/�hU>	":[�!_�3 ���V�Oq��J��C>��6�ͧc���ɔ�Rko�����յ��t�#	?,�*��a��uŏ��i��&�T%®����eǐ5��vApѕ�MC����r�z�]�J�+�_~��9��,�/\J�u�k��` ���V�MbOR�qAX:C�T���T�w���B�k�P�Ϸ��>��\uh*Xf�� 3�O��LY�o��P��W1���׉%:o�|�h$���5�aT�M/�i�#62��*�{T�o߯�k�,C$c Td&Z�	J��Xھn۫Q�����9U��M~gçb���i��;Vk_�Ŧ���Aۇ�-A����W?�� �M�z�[e���͖x�]����{���A7������(��d�e������eJԂ���V�ӑ`��ܲ�nq5ə�"��hMu�},iRHw9Qd���k����U�,����I��&)+|.f9S�*���
��
x��4��������x!COŽ��1loG�Xu�~Q9�w�Z~�hz�>��At`vk��~�X�����Ȏ4Y<s6a�Υn�B�]TWٮ@N݉�/�=2
9ѷ��?�X^N��߈��0����V3k�l*�Ѣ	h�%D��a�s����WZ�y��F��M$]Ġk��$ؤ��꥛p�[b	�R~ap���i��6~B�&%��4�[b �P�H� �n�m��%2~�EE1)Ϝ���&�⍌��c��ML�$�yA Ζ��d���ϋ�Ma&IC�x����h��%���X��	c(b�%q�$/8�HR���g�[���c6����Ŝ�q����vPQi����4.�`�֟@�S~��G:+�m9013��j����K���7ʯ@T �,$%TM�̅H"�M�C�����5��_��K�4�UZy�,�3'����8��|8�,J�0�GI_�������(��XӃa\A���-}�oq:����?���~iW��a�'���|��C%f[yIˉ�Z�A7v(B��G�=ڄ&����(,3$@��u[�﨨4�3�_�iM��:e>�8S�҄�3⳧99��K9�������ʞFe]��jֺ���"�׾}i�ήk.�\�dr<�O�a�i+0��Ik��m�)���T=�٦D��/��^��w願��q?��0j���P�����L��j���^����J��2�P��'�&��͹e��h�\>�'Ћ�X|z�-~���8�y��'�k�G��ژ��@"u�3��8/z�=x�C~9e�5�����Z�N���
��.jt���B7B;o��~u��'�?a,F�v$��N�f��ldfV7�} t���w$6�d�<�C?��<pi�Ĝ e�-^��6.N�	�?�}7�.�+���M�a�e���y
d0���]LO�B�<{'�X߸�`}�M6�]}���v���=�Q�	_����&��6�Uq���e*�ZNḚ77�Dg��F�n�:{�~�w�MhN48��T@܎&*����&�tdrdڑ���>�-�ƣ�p���rI|��uRV�+���*I˲~��22I	��9�y~~��|�ʭRQ�U�Em ��Y��Dc	e}����W�#��1�PmjW�e�ٶ�k�(9���8�,u-
�t�I����㽋8�1�J���.4:�lv�\�"D8j�=Y�j����8)L����H�=Zw��;~:)~dCk�ȴ�47�Ǚy�w���8L���E�}-rt2[B���!&5�HW�x3a�z^Jg�4�f��\���>5LTz�C��]�D��%o���^Q��)BiD���>����8���j���kk�7��8�$���h!���u����X)��A����ijL0B|]zD0m�7Ҍ���X*�����->����,"�0�T������4��[deF��x�[v�gh�xpŃ0a�Z��jʑ�e�CV%���Y��Ǳ4�"q�Ipܢ ���A��f���˧�t��g���j�;�/u=��(�ܴ�g���+���C�ja����+�[��"�w�KSJ}m�-�0g���)�&���ff�๞�6�`<|V�
/��ۣG�K`�[`�;w����1H?cnf���|~pwҩ���#ٺ��V77��eX�p�n�h#ZУ/�����ח�☊JV�uҾ�������)��Ѕ��a�Ӛ�̄\����.*n �"��M�V�k/f�AHz>�c��Um�̇���6�(�=˱�[_��^D2S/߻~��T#��IX��st�"�&FO}����j'f������]2���%}%he�,A^��v��1�Bs=����a�ţ����\]u�w��:o�)R�U%'鴍O*5`�h�tv���;��%�VŞ�|���-�84�x��������˕��=��<�Z�+���:z�6J�ҵ�����D� �E�mNxYڞ_�� 3�ymm�g�]���]Ae�z�����lL����@�/���%fZv
��:ϻ�wև�k��T �e��&t��43�^ͧ��7�*RC�Z=��L[�������$�3�e�o|靇kKuIEyI��ᆣ/��n�~QV���Mi�ӟۋ3@a?,?�"�cÎL��~~��#�1�*�u���_ҥ����T�����僋�V3G$��G<����oAu�	6�ap��z{���S�]�i�S_a�蕜Nu�"�MH�LIh��݆�V4�@NO�~f"�;�Y���g��T�&)�0�*�}�����ڣ��A����ŋ��I�m(i��ߋ����S����=qs5C��{$ѨX�-4`~�5�0���v)��\:?hukx�l�Mb���̸͈	ck`�
�=:�?������F�$sަ���Շ?��H�硈�Q���z�m�,}f�m�3�Y#3«It�}��n�4��EC����kI}��u��O��G��M\���w�i���5*�����,�����	�����v����;�زlH3���{f
m�J�^65����X��;!��C��/c&h_��t�9��7b$ �Z��@K��v�Y�Z��:�ge�)��FHB��~jʪ�7hJPD���L+Ptk��J��C$�q��NH���<T/7NR-��9Q�PA͔P9{L�:A}Fl��)cT#@�����=� ,����.�LT�������0��7�3k�o�:�1���D�h>�:/%��4[#$��&�ɜ�y�+!6�G��1y�3�*���{��Y���Ow�P>cϔ�[3���$|��9*�.������i5Ȼ��^ף�Sԗ�X�������� Z�(�u�n��.B����nz����)����P�O@�nA���.:�Aogve |�`�LꚎ4�bE�#���QL���8j�"gU�ЭC�U[��h o����	P7�0v|�\Ca��G-VNn�H��/h?/��}��ڿ�G2�]�3�$�0$P�{� *C�� M�p@�#��}Y-&��k$"���6���`�Afڍ�����')(\$�*���� �ρŎj�TiV2�O=���;���3�D7��%of�L"i�����K�~���r.t�W��C�z�DU}aI���>������.��ԐFޖ�������v�-�ޞK2��	l��^�{o�g1��n�Kf~�kW�r��#$b�z1I�6�x���Y�m}������<R���Q��/EmV(��8���_����j�bT�	|1Iu��N�����	q)�~�q���6SWH5OA󹶛hf}�F
7�*X���y�y��u�@d�j�ͣV�qV]Z�ݲP/�Q8t����)G���hVO:h#,`n�0�5�[��ǐQFE��la��+�[��KSbQ�P�S����� �;Pt���u�R� �_�#2^��i݀!�mK��0e����Ud$Y��I1Fj�>�K��Iđ��U�͑7˷Lٳg�Ѥ�ky,�
��\b�E�l���[�u����1�����bjG�ݠ5���^h��_���ĔY��)��gxB�/SE�_*h@*�>pp"ښ5l{c}/:��^�@���I�zơ`k��S �pNֱ5�S5!� 7i��ƫ�o�4�B��R����N+�M���#qO؏p�d7̫Iv�Xw4e�~*�P�8��H���9�Z	��ZZQ�YO2e�MXւQ/y���!֦}�#��~l����qv�4��'/��\��&����J$��xL��׊O��3�~q�^ugG�I�S��`K�'I
,:c���Kbi�[��iK�>ș���â�fQЁ>&��7�a�D
�e�q��l�)����Dw
j""eN���r���Yr��%`53���L����g���l�pBK�tS]Pv�u=���
�ĵ+)_���4w̦�^�T�T����%W���d Ui�,)I�3���V|��|^} ������S�ʋ.*q�9���)�o��M��%g�~U@kڙ/����P_e��>��~YM"�� :�Co�<('���pd���'���zQ������ծ��.��[C�FFB�N����(f�J4�
�i�F��I8ʶWgYg�R`B[����bFCxm��oX�n�A�-K���{/Ø�*�@��0!3Y|VK�n�<U���քo(�
����?�G7[0}��[��
�d�u�(�f��e�:/��#W�/�>����7Eet�I�k�8�Xy�4���W�[ݷo��җV
K����}�!;5,��)Td+���s�h�:%����?7�Iߏ(*f��s�f�:�{�����:W0��N5|�_O�QLx���j�K���"jj~�S�QW�@џѵ��t��F����xE�7��5��5�z�H8VE�GX���(�\�*�:��}vfS��w:`_x���$�z�u��f*��Z-qq����V�OS�x}���i�|�d���LRQaI��>��p�FkQ��`�U�N>�[.�'�@2�|_��_z���Z�(k`���~Y-����,�����������h�0��2Β7��0�viJ�*{͜�;uJ�'��0~�ӕ^�b~�68�\��_>(�S��G{��<5ܷ`�,��l�r�-�Ću��^����[k��gx%��"�-��#ش=��>�m�q鶜��U�O6b�"����%J/�w{q?�h=�'����du
�T��p�D�0h}��.���p��;] !Ͻ������g?����Rl�B��e$nb\�����`N����Q
=0�����z��呇����P.&��<k5���
�冩V�V���I��tC��ڹ���p�W�����h��&�..�~+���:'��=V}͠�WՎ߭��Q:l�6�^�	����[���m;s�<n.U� ��?=:XB~T���J ��\�k�t8\ZO�W�y�Ѕ�9,��H�>07�`��=���
���*��p��9�n��SY����-S��	��v(�t�����N��0���jJ��]T���<�a��PZN�
yԊ<�
��m�-�-iW��o{3���0G[���iG���[w��>���]�b�@��7r�b�U̭M�ElG���es�ȸ)䘏�I�����e",J��¼��^�)2?> �E��#���I��Y4��s-O=q��<�j��e��jL�M�3hFg9��-�J���}>vM	?��2a�S4�v�ֿ����mU�Q~"����}E��.Ų=�6E~_j��2�Mn&*��\���8șc��";Ѷ�*x���l�53� �8�![�1��f��}~�U?L�*��uī����aԘ�����54�4|�7��
�F�9[����w�P�H!�]�I������`��o|B��}W����̚򁲝���g'�f���f���ޔ����|�*�C.(ݦ$>�ّ{���S����z��
�`����Q#��B�����	�?���+;�@g�F<x=�&y����4>��&�U��"�(dN6E��3	=��yk;z�+�q�m{�6du6�v�G�R9�F�3��P�xe/�RC��xD^��:��-����9�0���v��Nf�S�5S
�*eݖ��K��N9�{.��/}0='�,�����E�b�>����$[z ������㷎KE?��Q�D$�CM�C !U>>��oh%�
�Dm޳GD&p >���>��q%;����m=�W�V#��Zx��1���?��(q��(�O���4A~@�G�b��:�8���W�t�P����O@d��CFUHa�h���/�QP�9�R���l�!��$��X#��	��,�)�)W7,�8-��s:��>�@����WFɄ�<h���rX!�����4��0��6"�#I����씉G��ĉ!"�#����q��F(ɭ��X���~��dx�pPw)��������u���>���������A���6k+�[6Qh��@�mO���oJn�'(`���nDa�w�¦���8����FM	��}J��X5]I� jV� :yF�\��Y�L	���őE>;T���DS��.d����l/��$�g������w����y�~@��EET�z����6��B�?�!��M�̠a�-��p�P����YE�9/*��e��<9Q�r�K �=��,{�ҝ�^�f�-�?X&�*���r��O���e{Q�$�  (��w���MpU�[���;~���ec�	9�:��v�6�'-	�X��q�B�_ChjC?h��-�R˪�(��xb,;���;�4X;p�n;O�x�+
yظG���ih���)�e��z!w`߮h��.u�l�I��į�ٔYf9��2@�db~iupf�0uZ��T��F"|%�ٕ�� _����Db�N��Hlz�}���'u�\q��Q��q�����K�HJ���B�\U����T��kO���'�\FAO<׵io�Y�����!�#���4��:v�:F��1%�;%�8����t�D/	7Jj��I�ƅ	O4��f�u1q��gA��wR@BcG�N8`\(�o����9�>k��b���L�T��V�J�4�A=j����_����[J�Զ,�}�3�[_�^�Z��Wj딾�1jk�F�]�Lf�C�`��d;b���Z �K ��|��L|��Sq^{�#�#��?Ȗ�_���=g:_�A�si�0���-��	��>��H�P'� ���g�c!�ՙ�ir_!��D������2vɟ��?�䟭�W��"���\��|OFu[ӥgA6�>����c[�{�#�&7���*���7�$��_%�V2K��X�d?��mkA5�"文�0��V._������(ȷi��S?"�P�[qc���;�KtY�U:JMc�}yQ�t||�}��w$��S���۵��a�&��a�c&�!hPo�h-���޻8S-�7?���w=Y�mΒE����ת�����ld��ۥ�p- �[�E#�9=>����7�8�;�9�U�yF��
���Q	QP����:�G9`*�P�4qv� U
�{�E�)z�� �ch	�;�z�צIA!�XYG	��H(�$��(��Pf��0��:w��ٛ��O�N�GE�"=���d�0�{? �+s���G���Ɩh��7%�?cc\ߜ5����
[Ǐ�h'}a�Ǝ8�E��9��2a��0�
��_��!$8t������p�ӈ�Ⱥ�A��O2�N��i��"<��?�(�q�8�E-�k��>hߑ|
�/�(?����;U�����&|+�c��,vv%I�2��DNlS��4�W#^`�̯�����Tg� �r8��U�ݝU�^���&�J=�^!R�4p�d�`#̈=W;Њ�19o>s��i�7�z8�Pq/��$���n7_N�E?� ��;������fc���օ5�{g�<#L�&J8Z*��)����Ϥ�j�����9gsIT��dZ_e�����۾@AwDs0,�4h\//�If���.��Q��L��i�Du����]8�I�
ɖ��9筈{�c�JqZ��Π>)�Ӗn�/~�qq,c⃚9{s�p��t!z
+�'���OIr�٭cT<���@H�"%̍�|��ۻ��ɪ���`�a�q�u�	�����n�����*�j;���ǭ� �ЍFl8�b�p�E��r���5��|��zTe��\ѯ�|�Q���:�!q��@�O��p`��� Ӌ���;��tr���4\!@��J�F�)�;0"������̾��5��+-v�=�w�ݍC89YR��$F�=�Ty|�+��S��.�����r��J�9*y�u�w�ں����U4P��ƬoB':��:r|�ћ㐽醰���*6-����UM%�B�!;��0jU�R��\��j��aD`��a�?x��B�������
	��hս�l��:��s��6:f���u |��.B�����~O��ەp����ʎ� �фHp
�"U��[ոt�t���۝H��B�%+������=��Ϥ�W����LY��~6�'�mR��f���":���c�DK=��]["��G���-j�}����RJ�x�ɀW%�כ�<1�P]��� _��"�K��F�l9_������
�����������a�B¯v��+x���!>��v5���+��c��/?5md�*RD#�*5��H;X�xfn^ec��[����n��W�7�z����aq�ŗWq�D76�F��je���N�Mc˶�8�:z�_@�[6�L�b����MZ5����E~�RM@Q�m7�8
w�h�@ Uo����|��,#7��د������a�����<x��7��*�k �Fib���t����v7Y\���  ֊�zB�`��'���\q%�����r���U��}�@2�Ҟ�����\C�)��u��5~�V����V��mZ}0.=b�����q 
�m%D\	*��z"òagƲ��:�|��N��o��at��F���̇���S��}�e��`?�"��źG�ǈAˆ���)�1FջD���]�n8z�y��YrI(��8��ǭ� }�uחy�[��C��J#j�� �}O���9Cd�)�u�3��䩖�
��������4e+�S�5����}-�^Sj!�V����1ͬg`�gחp��)���B�Q�A�xI��VA�w��.�K)4������q��� ����c���� b��+b����l��'��*�FUw�Sң�k&
��t�QD�o����M�Wg~�a�^�g�2J���z<-l�N���m��D�9��0H���n��yu	�ȫ�<��x�qĹ[<����֖�$՟����A�p�0��АܯI�� B "��x�����?�3�<��J��W,l߭�~���̗������*lDp��r��Ij�m�qt���3�0}�lЦӟ���l�v�����u}��l,�|P�e��*��|m��ZbM�f~x�%���%vU��E��Z��֐f	N��3$1d�Ɖ�[i�������cz����KN��i�!n�����iB�Q�r���#M��TT'���c�5x��'��V(����l���8�w�i��7�s��	pTh׊�쯁�~�j6r2�7N^]��:�����'_���F�t%Ro�.��,c	$ �U�Ԝ��Ũ< q?@hs�H���AJ&�߇�!��'�����z^��c�6�0�2ۘE�V�-Y�?4V3�X'd$����Zĉi�ƌu��f$aȭ$��~j-2Sj�8�D&>$��l�����������P��-�̒��T���LWx���\x��s&��5�>�y8ɥC�A�����D�&#u�KfѪ}#�H�9N1ջWG�Ә�k��8��2�&ӏ���>f<i�V<����I5;�糪§BV孚b5\1���t���D b��p���;SA�@V6Zr��*Q��ӏY�Yz�h��)2�k�'���eL�`~�U�)��KX�w*��
ˆO;%S�f�ҎU�%ꁃX���8g��8�^B�*E����y��C�WP;@�Գ~i'��y� (�&	M��ſt��.'��S@�Tx��Y�bCF� �B��{�(��D�#��L�(^��f.������N.7�/$`Y�����l}�y��ܪ>��M�n��o� �X�p��	Y��D.*w�1j�w�.�[�:N�P���{��9ꬂ����@~�J#���b�8�7���p����N�I��~�T�:�n��I�<�^o����$�����]��� ��7��Z\�n�lJ�d�<#�L7=L)Tv����
��������HC�_%�(�[]5�%p��5X�/a�����`Lj�`�/D8RN�*L�Ki����E�oA��!f�����-iO�s�i��I(��y�cE�Ԯp�&��'\X�0��V_.���I�A�x���fL�ȋ���-��=#}1hJ�i��p>eB���8�=d�{�In�2�w�l��0����
�ݥwj�"|������'|�T�;o+����X��iZ]<ƽ�"wߔ�w�Ol-'���$^�9	��9XG\)��G�"��֟szccU���ҳa�[��˸)��T���[������s�L�> O�$��=+�?b��T|�˅_H��=����h�������#��b�|���ҿSJ�Qve}��t(�='�x�3���5�kWZ~��*�M:��j`�W�r�9��|�e���>�-E��Q���y:�z?*R+c��3%�V�'�2��x*���]��"�5�\�T݌����.썾r�r��xm���f_{�'3�"�t^|���f�t ��=�zGqz�Y����:��Wg��B�U��&� �dKQ��S��V���@7�?��Vϻ���K�K�ƨW�{<�5���KD�ȍ�����1p�	4x��W8�}�a)z�\5���>#�6��ڮ�I��`�3RPOw�`?0��7��@PdR���Ӏ��~�Z�ٿ1��./���@�๺F�z���@r�C:(�δ�8�W���4����Jx	t��rMM�V ;���Y	��%|~�� ��?���bA�w�1{��S��-�ZNd�ۏ8��Z�)IF}c�Z�!�3V��l+w�{f�������;류�ι��~x�u�2^V�:=X�­����Q8Y���)�g�O&��Fm�B�5�n`0j�1�}�1��'�Ȝ�q��6�$��g��l���WѮ+!Y�5'0נ";���o��vU�}��9���k޴C����ʬ̧$b�=tJ}!�uCR�5�r=���4��p���D��̪�Wm��Z�;S9�o��?٠�ܵC�<fzw�1��7���eEu'�-�^�ݾ��)dc}��
rO��X�T���H�J:'��,����ɷ$�����VVI�J��WNͫ=��Ai��,U��	~�%&�n��Fx�f=�)X��k>蓷��O�
��۹�
�x1[����;�5r�%D6�<@�c�Χ�Ͼ�o�N�?�ů�+5#��v�w읰p�[������'5�����6o��Ĝ�TǦE�Ϟ���1P`��˴77ٲ=.P�R��ȃ��0Yz�� ��W�Ldb���|�j����m�h;hU����FW�0ꞧG���t��Q�Z�m�0I�S�{5ss�� �E���S�����Ƈ�$��߳A�3��{��qϊB���!��r,Q
�Z��	��/ښW��ɥ`J�쀓�Dv�駈����@
��ܷ�ֿ�P	R[���#-�������.G�d��`�ր�t���.�p����L��+Ԕ��>%�7?�1mZ 'y��! @��d��]�b��
���/���rc�J���w�~��������>��[����<�0��0��W�� �t�J�'@�"�>:.Z�Di���_��]܀OuvWl~zf�)~ʉ����6ߙO�g�kS|�E�ӢT���8��}d"�|��:n]w�V;+�2l([rS76z�0{Zfj ��!:D߸8�ҟc���`���9��v�9�m�VpD�ø����T��TS��iRd`6\) ̐~p��p�|wһ��𛝀uq��%��_k�����>+ƿ�nD/X
&ri��`�He�v�S|:���B���Q�_{b����-���,�g�9Q�{O�j���yz��K�e$���G�����_�gU^��@��bU��~X+4Ll����C#3�i�F�xi� ��Wn��p��c"Q�:&�S����q3H��+�ܨ��nCՍ���_+V:�V{�#�)��`/f:	�	[�tX%s�T�U���� F�(ߓ���$ᒭ�@�R
oKimb6�&�$U���@c�Y]:�Ј~�P)2�'�m	���T�j�T:lݼ�&�����]%��a��y7u@�X�s�2�hFg�=�1o0��1OJ$��0�3z��NJ����#�`������5U0v�ca�C�q�y��RK��[`��4W�W�
tep����f=N;��/�x@c�����z�7�����۰o2H��m�����Xey�`����?Y��A��HYW){<���!2�L��~ i�i	�8�%rQ@��W<Nn�-�3�	�IcCl���+�=�͜�V����t�~�0l��Q�d�3>�����͈vM����fu6ߐ��F�h���/0/6�Ё�+��Z�΃&IZ�)!\�2ct:��#ْ�qo�l�ؔ�� a��y0��e�����i��ȳhf�4,�ө�g�X!�Qc솒��J��լ}��L��{��������02�l�jCIl�fw1v*�Qˑp�u��a�>��`���)����V�7�ì����Bj�@65�l|�	�!�P>|���3���̒f�e����r�g��Ŏ�E���;+�Ʉ����=G�wcnI+j�w�	���n�Q�z"��7̇*^X��Sګǻ��$=����bc�<����ro
�6���e�>�Q�ѤP�Y�^�R��©;`'-�N�F|!~��rDNP?צ�
����B<�V��&�Z�[�M0�p8n�J��b<�Cڟ���>j��Q/8�
}|ԟ��� �E���D�;X�\	*�E���.�{s�9�C�ces�N8��]���ѭ��O�v51��cFG&X�CI�5U��p���Ύ-`_:������)׀WrToY7��F3�����od��J���<������SA����w���SBP��!G@�^p������2ۖ�~l�/@ylm$��=^F�PF���ư�7u��Gjl��{�L3�f�X9:��=�:*w�+�jG�fFI�u�`
_l�G|?v���C���h��L+\�<~�a�d�M�q����Epn��~Bji!	���F��/�Џ�r��nm(9н������*���u��+�|sPEd�s�=@ȷ�D8j�%��j�L,�d��D�u���k�F��`�&�*r��@�@e\Q�8�(V��>K��d�sZ������KZ(��Λ�]���XM�hu�dv�w\#3>�*^�1=�b7^�rb�x7%1�� s��S=@�	\$C#�u���,T��y�=
��2Qo��3���J>�B��|�*	E���r���9�c�+DQچcn���m5Xݝ���M��W�?���$��v��ZΜX���_ yb5��u���x1Ͷ�3�$�5$c���CB �j�K%���qZ�����:�mA���V7M~�Ȃ��`��~H�A����������d��������F$y��x�fͽ���ݻ=M������?1L �-�F�Z��L~��c<�CD���_XT[!h�bP����� 2�-��r���[C�puvsgr�;1��z��Bzv3��QH���KԔ��ϝ�Y>	�"m���'=�]��GO�YX���U����K>F��DuMغ���7�>Q}M�6� ��&^����o�����u�w�tS�Qj��$5��pÎI��r̃�ߏ�I�8hM>��N}zCK7�U-e��'���1=@�����f����xl���-�LGy��A��L����:�V�W��Nڮt�C�]$��>�^qYh*T���rx��=#��<���m���G�V�P�0e�ܶ�|
�,F��Jى�
K�{��x��7���xPAC���v�m�7�_'>�6��P0jڧ)��B�ל��h\}�ŝ��f\���a���Ķ�����#�S��Ć�5�t�h)K���+��<����Ĉ��(���d�K�9vs�؆*0�ɷ�����!9_�&d��c!���pS���}��n}D�F���f������n���i��Z��ӻ�S�J���ý���ǪRu�Y� ���f�{]Of�F�o��*�����:T�t ����	�gh�=$���t"&j��8���(!J�BR�'��La��J���'[b�m&f����u��-��FZg*���{�L�ff\�!x��W l�/��=P!�󥫿~�e�@솨�#��i/�.ϳ�E�_�mĆmHUI �N5��̶�8��;�6!x���Ě\��(X�����Z���a�����InH%o����۸�Q�Y�k�n/M{f_K.�p��r�a��|C�dV14���Џ�	�A�8�b��bsdYx��Aʇ5�m�l�? __~���I8����T��̺���5��w��b{��6�1F�;+����~��z>7��A�>�3g�z�%�o숦!�j���}	S������@��zLB�#!�9�GNo0P;Q��jdq:�{���L���pUy"4�r�nK���_fD�8n�W��vJ�o.����}��W�2h\;e\�mʓ�^1Y,L�g����ʐf�w(nB ���r����:���O�n�o|���|Ј���miG�]���ӦQCݠMF/ �Kf�y��A�SxQO~��j
|1ky0	���@x��e�IG�0�I5!^�@��3>pa�f��W�`��b�]�ek�AYpj�;%F��4J���JܨRL�|���2w�yP�:sCDb���1Q,�e���Z�K�K�h���\�������Mt���K��_
���Z�ڿ�~eu���#/%��K��%߽��E<|�����m�8��,jގ�nDmު����V�	�����|حX�����������@�L9�d�9��O�LC��%�)[|�17�5�~f(��ln�	��"�����Eع�M�t+��<����U��$���̑m���V
�{2r^$�2	L�يl�̈n�������͝�Ś(�^�A<~D\�wx�!S+��r6k��I�l��.=$vOPx좘�I���h��V��Iңt�t^�G"������ϚR4"�]8y���Rl�W�4���`�U0@9��T5tX�c;>�m�T؃��xN��y��q�.��&O������>�; 	�B�'��}W�IY��Fu~s@�ime��_�ⴺؚm!�+���
*�-�+-il{�MN$5+�Gf`3�(z?�� ̋�j W���Z�|�6�����_d�J(<��[r2|dYXd���?�>��/�*&e�*y���L��Q�U��[݌"�b�
��?P���_;L�J�5��_�^��JlC�$_v(�H��������6���L��Q��נhg�g#ƍF�AڹJ�q.|F�u�s��� -�"��F+;����3wٸ��/��t��afC6�f�|9��Ij b����/�5�Z�:he��)f���B��P�ެ��w�!�4�o|	[��?�.��O�����?(��S,�/�b�8F��>����';a�xЦ��%��b\+ٽ�l<<lHS���&�r0����(��(Ӱaj�b���W��7��B�$J��@x�;j�.�qs�z���]��:Zk�n��qI����Â#�Sb�*������)����9�SH�?��V).Zg�b����g�|�XUwr�q?�E;����}G��۵���8��Oj�x�{�J�s���l	��P�]�4y����)^�b��D,�r��w|KG�|�8��X�ND	^�"=#���x	Z̈�;*9fQ��VۚN������kާ�/ɛ?�����3f��)���bN!�"����Թ�&Y�i�0R�of���>.&��)�6��3�4.�������S�P��NF��_F�l�dW��
���B�Z�V�C��@4���a�gT�O��i DQ���S�1��,|c�ˠ���v�\�5!��%1Fsa�P\�~\�=�8~J�"���Lý1#���w<�{��(�]�Y�?��,�r�	o�'��,EN�x�r ����CT��I�"S�c�h|��K�<����̾��i�J�i�}1N7�J��l�١�HP�k��~��R�Jh��"o��;�R����$�Qx(2���?��Js�����X�J��cٝ,�~��C+�XP����,��Җ�@ �����V��E�ň�2�b��nj�s:*���p�<��ͧ�[A����f��fW����	�)��i-!��z�Ǯ� ���í՗�a�d�2�Q�"�|��{.�Z1���$Ld��'���_��j�H�gt�A˃Y���$ے-�;ϋ0�D#;�BD��U��1�-�ƑV{E����AMϰϾ����x6�k«i�=�@����͑D3S�������M�F�����{��Jm�ݕ�I1�����_䂝L�7�䐉܉�����HCc�	>r ����A����g���s2
����E�m��z�$��ciG����a���}'�l_�6���k3Ώ�\�&��ŵ�M!�����Q�WU�~5�1۞�e-N�����ȋ0t����:H~g��-�F+�*7�IKZ�M �xMjgJd��ۻ�e����a��Y $�6[��,C>5-t�I��;)���P�&�>���B>�yĂ�@0�Zm��OqN�5����m��*>���y��"{Ȳ���2.��	������M�0l�il�>\n�)'�v		i�V ���<��
��@j�[��%�,"-X��v��n˒$ �"��ڻq�� ]_T
�F���DGew�y�#}l�U4+66g_���W�7"d|=��g�g��ɰ#}�Ҫ>��m����!@�^ҁ2�i�%}�_4>|Q(2k�-�g6i�|/�W\;i]��L���R�,�x;�&�֨��|�	>zX�.ˋͱE>������|��&�a�f*B�.$�V�Z���hk�q�Tn�`<kj�4�<�d�M��\Hi1���0xϭ}OVj�{E�����o�ZLߪ�{�����)n���^	c�4�Q�`ǆv:�����&�^��~B�=�J�m�Q���"��с+��M!z���P�+u��eK�������x���WB+�M���ٗ0`B����z�;��^�eA�v��ͭ��cAߤ6�o��Y�Y|}U*�+U��e��>o�h��L� w!VՐκ�:��f����aX*/��2G�9:���I��ju8X:t��E�lFu
J�^����Cܾu{\-�Lܧ+t�L���X��3jcr� 	_O/_A��T0�^�Ε��0��Z:���K��O9*��%@ti8N�n!h�¥_$�2_�uF��b�m+e�8�����a"�s��R�8v�i����Y��!�%@a�ڮI|�XVes�'�>씲�>�=�ܒ��:�8��m�b��}{��F����9~dz_P�Q�k�N`�Bu������Ӂ�V�0w�b`N�(��Xr�i��Sq����G��G�/�~X���q��L������Ʌ�ˁ,���O`O�	�@�}��	]�z�t��h�U{U�)��@���\�nh���W����8r	1j_���t��q�r��K�\�4� ݚ�"�$�d�5���֤0�S��7���Ca����r!�݊	�Wn-4�_]�Y��lK����9ʾUm6˩�Q5r�(��d����43�m��b����H?�h�q884~�z;C�@�Ǻ�A Y� ��Z�jӢ�,B���ά�A�e�-��d�&�]K|��H���s�Bค��:�l��E�ٙ%�$<@'GOw#0%�a%�f�N�d�	�z���Y�w�����x�3� � �(�':��r �Tt��g���
"�(��r��s9��9N=�g�mc$�+��o�[��Һ��d�#�;_1L6�D���1��Fe�(Ā�sM���qf�3,	!���� i��ة~�.4������2x>ЗW忷y��V-���us��,�a��7y�+W�`+�C��Yg�k&�U.>�D�s;i�r��\T�D8o��ۯ����,H�0q#TJZ��c�<�`�Ҡ;y�7����3'���)�Nv��`ޡ���A%�y��9�HDF�ip�����
��F�SH@�X}�@�$�<ΏM	��E�d�{�'�	 r�c�ק,bM����c�|^�,�ӆ[}�R����4�D?�V����*-
����jˎ;�<���@�PYވ��  ���>��?n�����M[t�x�ј[N���X�ڜ�`�)�; ��|�g� �/w� �5��OR��5���O7k`�k%a?�4rS؂�)
���{ <G����=k����\(�TҺX��ɜc�c����i�^v왪W���!G&��:���| �Y�ARG>��r��[hQi��o8 �݃�"72��a����[�*�L�e��Gƿ������bjo����'�,T�wF�h�^��ۤ�ױ��N�F�I�Z��ՙ��lf��j�[gYޝ3��9�p�Y���:��!�n�y'�����"��E�X��R�x����aLyW�C�?!,�qA�\�t7*�$K��=	���0��ޅ�(���\-/��g���W1K�.��q_R�P�dη�ӳz{�˓F�<,]���R%�P�A���҂�=�P	8���ٕ��Bi��J���ܒ<�)��X�b�§���Y$<#<�-�Ex,����m2G��0z���x��_��~����� �o�1�����(��Ϣ�� |�O>���c�ՠ���>(�������]l|t�<q��3n�����y����6����R�i5QS�.�'�Ɏy-4k�e,�-
������T�y�����3�c�M�x{�����h*/����Y`��tW"�'���<U�p�\�L.�]�������{j$>B�u*��C�����*k6�y�}���(�b�֘���a�Jt}��>��U,(�@> j�&����\�:;�YÛJ|��ʓ��0JL�B�[�A��;��A�5�%M�q2���: ]�J�VA0�t�#I��g���գ")F�0�&�t�\AvB�����8o�u� ��Kt�R	w�����(�@�K��^��|:z�Q�����F�>i��LD5o�^|�G7����U�줻&RYn���EWg6رaԀƹhx������^hR?�U�I|0��	�nT@:�v�=�~ �#��hc�Ҝ�;�{��\ߕ��O�+LV�U�uJ�"Sc�1���}�6s21�2��Z��z�4/��6_F��k���iyN|ÔW�z�i����^������T�X���G�x"���E+;z>yϾD�Ⱥ���!F����	���m.f��B�0�p>O�k5Ln�������Ye|\��L�G;�<���sw�����%�T�����/����Jz:;��:Vj������Es�V�=>C�dV\���y�'u�s��N{����,cz5�{�Ѹr����U�c!��O���Rm9�SC�������Xl�l�h.Dh�B��mP��E���~lE�A�,�8��F�l�\�������\�>E4�<�x��c�Y�b�M_U�o�f���H��u���?}I�s+ΔkA3a�'�3e3�q`���{m;�4��1%i络TL<�j�/d���X@_��v�Y�ß� #��`u�H�[��d�A�����x4�5n����vu���M���I���;O'�诡�6E�4$�i���6D�9�y�����1��1ct���vE�H�
YLyM3Tl�����mzo�/ճO��3�A��-(���U@��
r�I��r����I��?�(6]�j��Ti�Z�8�!�o=:��O�d���D�a��ö ��>Ź���{���V�]|�!sF>�O��Y��и�WV��OW5O���q���)�	�BbfaO@i��,��&�a��g��q��ȋf���њ����ߎ�Qy/[���N!�7>�~��� /ΤnZFop1�].@Zu��v`Y��|�w�jml���`k���
�e*'�ǜ�Fsl
'a�k
�$��(��}E� ep���9L�O\
�3έ�Hb�g0(���x��],�"���;*V⁃"��zAM�#1����6�<���H�RB?�q+a��z��Lq�H���z���>��S��-e]�b��������Ў��`���6�R^�ڳ�Ak\��)2ÂsJ\��H�=M��Ê-Ê���Fӫ������cq{�F��o9}�"TM �7\�_�èZ�
�g� <�,z�i�l����ڰ���%�֞L��m���*���i�Q��d'��Y_N=`ڊ���$�de�^�*���I��&u�ʠ&�U�x�F=����������"�`�Ū&N��7W�Z���j�`���lEl�l����w��%�x[n�u�R�kU���c�XJb�� ���=;�k���6黌��{�Zk<�F���O�.a�W������^}���\*烹�MB����������j-d�����N;åw*t�{�mrDrS�#&��d���V��e�ݑ��35/�I�>,��.�Z@�a��������bw����<���~H��-�el,E�^(�<����@�1?���S2��iS�ǈ	����O����t�����(Vgc�R뚩��x���D��5ia�v��'�@a��@MkU7O���g�K琛���o.� �|4�S<�s�nmd!�l�[� �<����7cU��R���+7�5.�Fc��'�uA�k|��b�4����>��5r(Df�� ��I�������g$*���{9��V��~����/?����_GT������K��ݕ��� �t��Cdzr�j3%�zP�	���&s<�%�����	;���͞�L�T����8#܄;K�e,D���L�Wb9�x��)�LP����`�(�s�n���X1
��J��f̂��h��8IF׸΢u{$��d��k ��ڵ3~%��%�1�ԓ�p�S�?�A����U��c�n'�ЕX���Kg�� �%yJ�Ū�I�g�|R����/E�+d��pc�^	�5����b�*�����/�'�6랩�ZzOx�XІ���� �/⿅����?������5���"?�.����K��ԟ'�F�'2v�:�Lo��Xe�挕�C{Rg�b$�$������W�9��`����;��-[��ï"j��b�Ӝ�t����`�� ���܇��� o��Y��%"�7'8��Q��N2��ǫ���.�����y.�m�V{��gi46ܓ��t$?בYMҊ���o'7�5��T�Y+S��)���J�k��#�����������zՂs�"j[9��5b�x��˲�����N���o��i)|2R0?Me�o��s��R% ��F���Ȅg�'h�`O'�;j��c4f�<zo�	uFm�� o�Q�kx�����eJt0�8��ڽ/l欨ё�2pY����%�F�<f��za�8�/����R��.��;8E��P��b�{�8,�	���/LS˯�]@�z��	���O�#�Y���d�����j�a��#���O�t�ilқ����9��Y�U���#3;Z0�	��a��T���Y~6~�ӳ�I�z=a��D��)�@Q��	5)m���4{�����o�!yz�����ڸ��I�q�[|��(	;��/�_�G��H�ˀ�\rN|(@e��s��|���^���[U��b����7�ͩ���w�o�ϳM&����Kw�F�{������cF뜊 U�X2 "h�-L�;���!Zž��S�};?�\qʈ����^P�c�͵t�A<��/MGv���M�ʹ#�����c�*��^m��1M;$�t�����������J�ߵGP�k�� �R�:R3�b���9�@�þ�%b]��N2@Y��b '��D�_DQb���n�����Cp�Y�u_��x�o�ŴF<	ux^��4^���J����}?�)UT�z�%�H#���& g>o�օ���˔���U�}�$��J�ܦ����+
�cA�%p1��!)�[������o���"�z��&�L�e_�Pd�$��}�8�������a������$A����yI	�$=�&@��b�=T��E�O�F��K�R�����1���΢�i�Za�����\��O�⼗[��郺Ib�lZB���l�0��Z�}��O>-���Y�it��y��{a�P?�Z$3�C:��-K%yĪ
~wֻ�U滑��)낈ez���E.B�aPusp$W�"��Zd;Kf�SY�he�kV�5FD8�B]Ns�6�'�I�d"����cK=���֘�m��n��m3|ƅ��+'�]�����uj(%�!V�}@ru�ku;jn�7jH�Z,�'Ia�k���L��J<� �B�m�W�g�ǡ]�P�%6N�)vh�_#r�E�%������s���K�`P�d��(���6���$%��Qa��,�eg�]�!3i�*',`w���b7nMH���X��(ʯO�4�Gѿ#L`����g̣�"�W�v�%��3�����?���YQ�H�DD�4��*U��3��K/I	yr]��W;�d���K3!t)Ö�h� ���`�ݰ�\QMj3�g%�#�4���x��*���������EO +&	�����g����`IL �2���&esw��3h��΀O���>��$�c�� �eq���f�YJS~c]l�g�ħ���Iv�zF^2Y�h�y�
hwXOy��p�J�մ�;Zi�_]G&����,�p���/~>,��L|����׹���V7$�$Uz[���Y/�ޕ+F4�'w2M�4?�@>�RMX_$h�(��X_��L�y��j�H�z>��}g�]�)���dަnX�~L���<9і쉏�e,\:\�ęY�	X�D�
O�@V-���}�xք������Ё�����ˀ��b��3��hx��i��ό��o-����K���26V}@F�����#v��Eꋡ㓫��%=-�J4F
0j�k�FRT��i^4�s8J�Ǚ%�B�@��������w~�����<�� ��׈�a��"~3#ƄI�,4q a��ц=0�/5K�ҥ��P77�,us�Q���K��o���%����W��)o�*QI�o��d�Rh�\(Ӭ������K�dB��B�;�����$�[x��{���R2���Hu�]o[G�Etܷ�$���f���a=��K�jKy5��-noF;������l"%^W�_a|�̖��IG�:��U掗�5+��n�+Bo6S_�����-ԼLk��4�@Lu��õ�b���o�cO�i!�L���aM�F�����c��Q�#��'f�����PSɔ���uB;���O�����D�/�ȿ@�0�K���=DDq�oF��C��D4Y�88խ�7!������c���g�3�b�w�gM|�K2�ʄ�˸5U��sH���C���@�@y�뙎m*����魝b��c���k�u%�oaE]�[�8�J$쀥9�.,�uz�G��������X�ٗ����<j�o�!�r������F]o�%����.ʄ�$�m�CY�A%֕����j�8�[98�Ka{���<�(�������6�p�XS�q.^)>Ȑ��X�Mq�c����;дu^}z�y#GuJW�����2~=y+���"��N�q����
_�tFR{�FD,7�����&��k����d'tW	�2�.iv��
.�^9̡�"��J)�*$��OD]¤-�Fv�W�Z%P�f#	���s���D3����!W[�.��_�E�	�e�܀�{tY�hWӾ8 �sm"�kP��i�H����{�Y��0Gf�P��E�����N�b v��|'�Pj��r��~�����h�(���}ݶ'�U�mɲю�ڳf�,���C]���$ն��n��mT���� 8S,��8d�q����ŕ�i�~5(���^�t�)$L����C�}���+&�}{\$ˎ����{��4�#�s�1ٚ�hE�W�*�ؤ-�Xw���FӢ�̧�S�L�s�)�qRJ�g{� �4���Q�8PN@zmۻ�g��m��cx�Y�c/��5&^}t0�5�%/��Ғu�l�a'`���΍`l�$N8�64�u�|#�jk>�(a��m�-\�&I�jZ��S��fY������W���(�y�E3����z�~�W�����)sW���μt?˛8X�qt�w�۝�g�?���#���4WNrjlq�K
�ح�T8��3�`�S)����ٜ��9ע�1�hsL�N�J��
@J8�2ߖ�u�r_S���&CW������R���?U���@;��`�}}�Q�F�����v
g��q�g�IM&��i3;:fWK��2.�.w��R9'}b���/8Wy.C!�������2w�Wa���z\��}��j�+\߹N�VqB.�S?&X2���~M�{��g���3L$��h�h�B�o��)%����s�8K�f�ս*��7�\7-K��
V�(���4L~�###�a��,��"�{E�;�]�^��D���?2�͂`X��ݩ��&�!�M�6�eZ�D����8�=�̺+���x�%`�D�w<��<����/��J�odNsK�XC�kbF�\�F��j� 0Ǻ���
@�q;��t�Z�g�%ym`�/ Պ���Cow����hɌO�V� �iF3�;���H8c1�fTW����e�)qp�伍{���I�~���;\�m8 /�F���{�/�CD�&�r-?g�+���
��f[��i,��/���H��ih�O����W��y`����[*�=�Ӊo����S(�kX�xuP KS�Օ�mC;�c�:���Wܚ������¢;�'sG/�K�E(<h��N�M�n�v�T�'� -�9�$�P���:J}?��+�PAp�@��̏g��|^aפ��l��a��E��D��
�qn��X�Sk{?uG�߸�wz���쏁�oY-��m{���B�8	��~C�15�*�#{���%�Z�7i�T��B�#J��W5��G\Φ�r�ˡ���A�3�^�1�%Z�ٺ��w$r~n�0ǈ�/i�gi>��r���+{tW�U�R�(����Մ߀��#/�H�p�Pn���Ȟh�,�C�{�>���	��h-'��I>����HIa���cF=$�L�y!�K
m�Ne��gxJ�x ɲ(��w��>�C��La�ִWb�Yӽ�Y���D5<�hǍo�y+��l^� ˯�����?Z'�f�j��u $��8�-�.��e�ݤI����`�ӯ3F�v�Z� ��d-�~e��!�|\�URm�t�]�6��;p㰉-%��^C����ш�9�{�C�`�%\��K�j�\������ X���:�l39rR�?�~����00A������!;��I�z�^y��%�܇EZ���C��vr�n��@̠�&&;�,��G�Hp�[d򤻧�(���k|\�)���C�G0�3�O��K�-�� $ ����H�����U�l��Q��B�4b@��0��VX��i�v�{����âScyw�e���OT�%�9�"&�����<�sr�d�H��Rҳzw5}F^���BZ:=��I�������'�ܭ�y���i�+��z��F8Ƴy��
a�o5�im�nȲ�Z�s��`� ��f��y�rkSn����>��RX�X��%��>�/��ڳ�B]�����U/����^%�k��(�
K��� 0%�`�
H*�:�b���z�WV��j�f�������/�j���ђf�:�EO�eA�)������h"w������|�U��F���,^~l�H��s�0��P0�-�3�q,Rd�/��w�h�َ��(7l�?èr}J�-��-vL�>�MfR;����8��o��(n,���kqw�������4�v{i��=7��Y'1]ľ#P/�<,/[�uS*��+���1l �� EG����`�B�f�퍨�X��*�ލj��l�Tnf�\2����BpG3���8ȥz��S�<g�r�e�[f|n�a��N�j�Ϸ�F��C*��rT4��C��R`��O��r��F��a����q�(��x}?��I�� 0 dB6w�aFЋW�?<)
�R�\[	�l>�:�S�pF�
Kqؐ��oK���خ��Q�j��fˠP��� 53�5��-Ԅ�]lT��~Ǡ|���V��a5o�k9U�gQ��d��,0�c%8*i�	|F0$3��}� �l��̼�J�'9���%�GV��������&y`���=�S�s|�/s���`��7TA�'�ۈ��[�u����{ɞ�)�QU���E�C��4�+O�|:�ڎ;gk\� >{��7A��-��o��J���;߳�~W"��:>�SF�l�y�Q#x�o�g�����o�?�D
���%���(o&x��/�����^��JV�$��im��Ȧ��9�Z��t.�'C,*)��o����c�����"u6�|�!n�R�<�t8�$m0|\K�ՠ�C��|����@���vd�3�լK<����PR��/|Q��P*�6x۪��iK���N��N��\�,��K`�9�f�O��˼��~T�0�ɇ�;?A��/�^�rȥOT�t|ǔ�Yk�Ĺ">lT�M)gՖQN��F�^�)�X��0;����	�t^BN�&}������]�=���N��K��'� 9J��[���c_��e��3�n��`0e���$^�w���B7Ca��S��r@�Qh�t��o��r��JBt�9S�ş,���1H>��ch1z�4)y�)��u`?�X���#E��b�ju�e�^��P�������: �]KZ��DQ:1��l�=o7�8��1 ��!٬�B��LEF�r�0L�'��Y|-�e��EG8|u4r�AYO>F��#$��다p�������M��6^�ym�+i���uU��i��'�b��V�VU�WR�BSn����zYH�C)f�I�ܻl#��p���h?��dG�S�/��wEI��eHD>��ퟎ�2o�6T��45�4#��銸�w<5�ʸ�@�6b\;i_�!�T�<�U�7��e�S���i��8F����N[�U�K.G�9MQ}�|����Y���JՑ=&�8��p�3��h���"�F�T� �s!���Z�����WA�AmE�"�L՛���A�dm�
���6��e�y�QP?5�;����]a\^�2՚;�_��uW�O�j/��A���]'�Ϡ ]�����"��;��[���ť�K��0� ���|) �G2�&�rqw�f���=r):Z~�� �'�
��r���g�>O�#0Z©�Q�&�<N�P��P���l9Z�?���D	��?����A^E��PM"��?���է3�{PD�Yۜ�]�u�?A�R>�Ԕ&����EH�VL�<�{
m#:��|,l_�������9���D4/�e��w�9ʯj���<"oz����#Y1��ૻ�Yu`y�}����eՍ!���hl��5F�7��D�j]��[�sG)�O�|��({�[K{ Ƅ_�Px�s���@@����I�x9����k�=��q﹆eN�t�k�(y�C�f{:���?nE�����B���Δ?ߝZ�-h��	ԓ=�m���s�bt�����[y�s<ۢ�W���NˈQ:�fF���	��^n_Sj+f�&���bk����#Y"��ԗ�DC��T@���2:�=�!��mѐŲS�������;^*��!_�
3љL��H���������j����ֽ��s����]3P�ׂ��]�N�ܠ+s��s��j?�pč��?�-���ٽ��ԡ۔���n����u�{7����c�+���gh��o�V��u�������N�� �	���*��8Q����`eD��wG���C��ľ ��n���t[���g���̋צ�/��6��q��O@�Y�7��49��8{�pg%L�}!��P,G��.�Z.��o�s_�VL�_����%��M4Oǟw�n�z�;���O�1X)g��1~W/��������<P��T���9Y��JuS����� |���*��-����Y���j���=v�������_+�+����tc��*��O]i-f#T��W,<7D��#��)��d	hP���1K��IY����r���A�P2�;-����O"�����=����2� ��nPx8r�_��(4���(R�����@I�pF�*��5��H�sZ'�r-j)Tkx��p����+���g��i��n�
����;�L����1��]_v�����uH���y&��wlh^��#3����xS��<�O����:e��Z_�at9�f�q��N���0�4w�|�/o�H`"�a���O���S�<�"\��	�U�\��'X�&��f��G�o��K2�y�/�Vи-��ņ�Q��z�L�u��g>���D�*�K��+NYjS������B�踲�weu�j�>��7���y�wL���e�o!��p�����Xp���i�׹�lXH<�chz���[t���Nd�!�����<+�S�2XMʜ|*b;}Z�E��/-����׏���F���'x}?��B���6ɟ�:d3$�k_�����<���Fg��L/��Y?�8�������ԯS��Оn^G��U �d�m����343#��x#�L�}H��dw ����H7�Z=���?e
]��FX���7TLˏX��i�G���0�K�$�\���-��s���QE�S�l"<0���=�^����k�W�PY(�M�����Q�ҏ��_�����Ĵ2hz��O�b��uq���l[�ܼC�y��eM״���1��B]�RmS6�Q֓��m[�s!c��D�<�d^�T|NF �l�^���~H���-�s�0�nv�o�.0��Z\&X��|~�	}+�<�Q��׳����Z�	���ơ��v5�ǐ�� ��7��rחvʂm<� �U�͉��U���۠JS�ۣ�|���%����'�p��}��@�Aۼ��s義F�/�m:�7ndG�ۙ&�\�Yz;ȶ�j��k�j������G�X2B��fc���h�0]qH���J��H���b=���@�0�k�q�>�A��&�t��ՋD�vn�Q��࢟QA������4�R��ï�@fܧ�=}4�l����'uӁW�%�3���].O�6-���u����,Ԕ�f���!�,RY<Mz�9)?�^����ä�G�����$����G;��U��J����դ��R�jJ�>�� ��xR��$�bJh8 '{c��#��B<�csN5
.�500���T��Xǯ"FJkY��k�Od>{�pz���^���M�V��l8��D���W�&�����~z�܏+�JUщ�8�˝�Ӻ/[��?P�p��cNm�TV�dCM�������nk��!@�"=���2ܢ�L
����u��(��������=渖 �d�W,��s쵀�r��%5<������7u3XM�ꋎy	�L�������%�%|x�R�jgK9)I�o����7$h��c)����6Vz�
��2�l���cyK��]9�F�F�}2T���s���(t,��0`���P��um/�`��x_ik S~��Ų�(��������鴉Q�}'��Gι�ɵ�x[cV����s(������5��t���;|:� ����2*�J)���r��Cݼ\�v�!���.c�р���K^'�����ϔ����w���!1�7�ҋ·�[٨�;!Z�qWoJ�"Y��1ba�U�)5�+&�Ƭx��3<�醂�f��1��͈A��Qӯ�M��}I�~�fs����9#���r�۹�Y��<4����B��+O�sr�3�Jڞ�J��g�r�l��%. xn��4Ƃ�<	/*��Y;mG>��U�3.��������c��s�����2:�א�ɆU���4���)�	�χ�)�<}@��T\$��'[5xR��+���?���[���z2a|�󬿭�,t�䎱��j�І&�s��m� j��W��K�sjhZG|�(&�b�u��K��U4��x�L@瑂��r�sJ�[8��+T2y�^��_�f��Bo�dc	r�요*U[r�<{�R��	��%��%���v�?/A�����5�9۪�OK����k�L<�$�Y�J��iU	��W5�L�q��i�9%#y�y�j�PU)�	�����Zϻ:X�v��x�o�;>o)R$J*qa�l<���S����I�3�#b�3��K-6�����ln�NP��dB3�៖b��h]����c��cKIԜ���	�7h��I����1Xr�4��p0YZ�?kŏ%������]CC�)��_7�:%=���l��7.ٶ�X�L�m��G�Gl���*}`��h/���/��7�i��()�����e
�T`��r�z�tώE�\�UCA��j�,	��.�>�}�

;�=7g����k��#*�N�W�:��mi��q6R6#
@����m�`��z�o�4o���z�K&���*�MAKabNݒ�kh��m�f�@K۴+��R
E��g�f�k�����gV"�Sܗs`g���b���]'��k���<���$���ՆG�N_��*�Sg��op�q� �GU�qi��e&$� AG����@E�#�hn
h��������j�f�֝0��2{饋���X�	��!TX~y�d��ɖs��'W�)Y�0�d������FK��u����La���&Ȉ��d.�S��r/�mrLM�b�ᓕ�+�}��͇^?j�,6ժ�U�C�o����;�;?R�7bH��n;6�&O�����}�^��	z�k�q�)B�����)j��e�on0D�y�{k��8�ܚ���M�g�6m�R�%6&��P�r�9\����5{�|��Ѕ�n�[~�~f��O͚�JI<�U����j������Зh�>$�ƺ�3,xtpzXx�
�i�L{������"K'�,��`��J���WA�x���#%��!g�2��N}��iψ�gGK�OA.�K����L�,��n�t��,|"�!P��	b�|������p����U}D�� H���b�t��v�%%���|@�9p1*~]7����
�*	,���:�,!Np ���3���ʾI�VM���p�"q���T1;��]�v��,�����t"_�*{�b�s�8ܗ~Wԝ�v�ޢՋ�� u
C-����'��){����]� v�Wr~�,�g��!�\��%m����*�ޣ=�����L��~�J�������#~AK��p�"*����o���ӛ����^�`��綧����lG�4tВ����ׯ��Pv�Ƙ��J[��d�<z�"�����3�N�9��7�C�u��I���u�toH��O�[��`�S\2~���?�+:��2��ޡ�@(5�;��B^G��Z���MNr�E	T�{�����Yc�*���c�x�s.�\D)���׎����A��r]+
��0�=#�J�tuN�t���2Y�jԎ���&�6S-���p��LX\;��Et�PYcmC��2�N\��ӷ��S�`�y�>�u��(��V��ѽ:�jd8�v([��%�U��?^V-�-B������1~�Zj�������O����O,]�@xnV�O�q|��7���	?�͢ڧ��88�Ļ�� +]-_��G�
zw� ��A
�}u<�"�;�R5:N��E��Y}ݔ�%zH�a�)��0;�(�'��ku6�~C��f3��Hu"$K։�����xcE���;�j
*�k���y ���:��o�lB��^u*�xM)���]���$u��yK��/�	�B����O�����n$'�������3��D�52Y
�u͏��H�zG\+y�����
��:�{e��n���V��e�p�D�$�q�/��D���򜂼�p�>Q�f}�H8�Op�����W��a��"/J��|�X��HL�p��o�rP��°	"|�c	�soA
렓�qIV6 �b��UG��A��}[�0��wK�v ]����OM�,L�����3q3G�C�"����M�1`�X�p
���Aa�2۟t��e�l�+��7��A1��m<N��$η�K!�!(%���k������l�%�Vjy�=d��c��#�@>0@L=e)eؠT������3����z���rƣ!Y��V�R쩏~��NOkAPc�g�k��[�'�Yn׭��Ifk�>�C��Y �\��[�ڎp�t?]������v+��]��~#�p�2`�9��:����^�mZ�7��}U�g��<>H���V�۫3�v/_"��zBG�} ;������혃O�he���(J�"�0:;|P ���e��� �MM�kUwî�u��/��z�jA�����* ��ɪ+�Æ��� CwѪ:oK����:'��!��L����m�-�VC(t�C�W�ʗ���7%��j�5dh�Ut��^�pk@����J����� sv�3c��i�0�m�컾*,����Nzb�Rq�\�~��O�c���xRY̳G�p���gU�a�����SωtI�"�KK�oI�'�џo�x"1lZ=%-����a���pM�2���g��Jײٷ�}s�U����CHH�.��b��GH͑)���� ����h�X�&�	m�,)8�ATk6�j�d��AA���Y��14P��r�el���X;f����	�!��^V�����H��2���(�]��~���D?H�@38j�9���҇��5aFMRf�SR�y� 7�%�; ㎱�)���eʑ�f�c���Ibw-'�[�q-Ci�Y|n��pԩ��c�z���H�TH%�T�ծ���%s����1H��@࠸���Ӯ �!p���˜�6�G�o��r���(J 5L̂7@�,:�����)V~Q� =��Csfa��ȂyNW�|ǈ��C�B>��D���k��o��z�>9�`(E&�(ۊ������i�l�P�5Ռb0�����3�É-Y|����i�����6І�G�Un~�@���kHv?��!qS6�7'��(���ba�a���7�3�zD
���%7W�p$���@�n)>�f&M�?�P�BD�'�^���gx�������N�&�e���E)%jp�����ξ_]��Y�(���2�d�T���!И���3z[�.�6� ��6�����.?nN��BBy�x!h������K�����;���R��3�ZqRL.,��P���c�gd4te�t�L��r���Zy�WDr,5_ ]h\Y���G�%�ݏ ��W�F?��d�,�o�X��j�N>�+n�5�F��k�L�h�0�LZ__J���qҐ�5m:z��s�NP8w��fNh|� I��k���ʞY���83�F'���\0�مxA�=Do_J�Ֆr���ߢ]�ܩ򒪨�U"�#�����1���a���7H$��au�n��7���6*��&_��u̝���U�|Lк�EY\	e�ȭ�7��˚�#�%��4�(|EN˅��3Nbc6�p/Z�<���%?����^����[YX��fP�-(��~1\c�G�r�\�����8�G���|�@���䀘~���3%���Jkiy�ð���'�K*+u���"�����[��<�)���7��U��Q_��s�������Ŝ<���� ��Rc�	�X����G��I/�ӊ�ax�k��l�Y:А*$�n��f�볽�1��	.`b�Z)�U0.�����h�t���IR:��1�F��w��+_/1���M�;���yW�a��R>ߡ��6QM� �ƜK��)Ӯ�Koq_�h5�N?�<�K�b�	Ε+Z1ne�	 C���۰�^�bЙ��E|F��2+�J��L�wiF]��թ�����H������NS���b�o��08)��!��a��d�"��u����
�(C�w<�(8���~�hݜF��ղ�e��ąV��wQй�8<'��z�}����]J��T1�DS�_8U�W?Jw/��r���$�5a��=�Ș�v6�G��	&+�cc�EЯ��r�q�[RT ��D�g�u���t#�c���n�9�P���-�/���e���g��f҉9�����v��¤Θh�Cک�����4����X��E>&'Y�U!��:�c+�=a!�뾧��o�Q��F���m`|&+�ﲿ������H� o�n��W��Y�큧�	I��.��7��%�%`�z)V07<�#��,7��|��������s�Ԑp�����
|a8�/2�B�eh���<�=�{i2��ʋH�p]��,ju���
Dn�vgB�:u?߯�N�R����Ll�6�3��f�2�/��\*vT�3�""�2"��m��+�sv��)��H�G�bcuqbe^��C�J
���b?͞�GHrPg~JX�y5�����K2���ge���-��Q_i�yqNs����Y�e(����"��%����dH){T����WSo����^�gP���j8 ���|`:M=�,7|]\���6�w��[���������1aĆs�ePDY�����9�+2G%���ʋoI$6w�t��{�F���#�t�
�U�_Z7�G5)5�,�B�IU��>������`�s�v��};�U& �v�W�j�蚣��q���>Hr+����su�_�UR <�w5��{�l0�����Ҡ���s��R�^�6�C�r����xuӭ��M�<���\���F��a������ь+n�c�QfOr����-/oK����,Пj��V�ۣo�d4��[bk��l����[��!j0v#	��=�O����L098��P1���`�Qx&1�Cu�Gl���^� ��M�/=L�^�ߨ�4�C�zu��1�l��� x�-��|�"����m!'��i��>���W��	��SWI4�&�U���93��r���4%Vn�����@=�4RocF�l� �{li�-��������H4��	�%,�m��<p��s�%�wk�%��ǌ�r�xF�,�+E��/��04����)b�^rl6�s��fq6t	Rj�%T|�����[��)Ђډ���R�=v�:H�<GpU�����EG��?�g&)<cYy���AF�w�rX��nH��]&��8?[��ی���ke�ϴ���_ËI9} �j%��`<F8K��ϓ�M~)�2(6]e�f-���?&�������z��YS={���Y�Lh�x��+�K�c�>�u�����!��V�y���^��*7�ч���8_TF��R>,cJ��_�;�Ԯ�D ��kz?��x�hkL�0��ʯ��}�j��5^�5"����"(���KC˾1+����ߕ����b*e�^��>@�Ԭ�(�X��.,#ᙑ�k�l|C�`v��&�;�Kf���;�����D7�x��ݷ}�nY?5ݓ��o��~���� ���ȍ�z�pZ�v��6�1��Ʃ��`�6�)%��M������^��0��B YQ +���~�]�����5w���Q����N@�w�Xǩ����	�}�ϲ�[�٭�-����)�ӃR�UH��o���뽝H�6l}�>�>z���^�fe�<�9t�2HB8�8�l����S.��}=єT"gʩ����	Qƾg7�0���g�6��}�������L���� Gv�L��u�h.�m1�'Au�4�C���n�n7 1�3�� �����ʐ^��5+#���j ���a6w;���^3�����|F`W�Vܪ
��mv���\ls�u�0���f���G������.��%�oi�H�R��$�4�c�����#��A�$�;�b65F%T��z� t�83�1�g����G�$�ѐ�܏Hv�&-�FFJ�w�w3�$eL}^�A�����s=����s���5EhR{5��Ŝ!a��&p0���R2��������ij����0y�w2�܃ ���p�/c��x �����YN�lo�{���i�4�R�߈
�)N7+������E��b��PdRYm�r�vmѩ-�+R��a�5L�-A[�0�E�̙�q1Pr�%�j����Ax�"v���j�i�����(GPKWx��0~�y�3g�I�}"��P�hF�.���@U�!R��	�,o��c1y�/����TH,u��1Գ&N�/z����������f� ����䗋��j�DPJ���/n��Ώ�4|5#�6[�{��U�R͐R�[4�z-`���j�X�5�]j�`5�Z$�\!�#o���̮�9E�6�=P ���*xsZ�M���Ԑ�U�]}�}�^Q9�!�Y�Tι|yր�;H�4Z- A�x۫����<�2��l/m��F�Q����W��	E��[XHl�PU���L�Z��\x��̍���OV,p�_:�TI����?]�uT�Ub^Jo.�Ax")�r��9j�$�4�ԌN��6�k�a	���T1�%ɵ8v���m�-����������K�uVzH������%@�ų*D�}�a{���� �N���Jc+8Ԝ���?�-|�X�H�'�Q�q�7r�h�j��^YqW:�i ����*R�vC����f<w:��mz�����[0���C�R�&mB#;u�.����@+������S�TC�)�p�(�aaԡ�%��&�X��LL����%�S�pX�Btc!�/�Mʋ��@O�+�x�S{��9Ul�P7��䝗߾�I��RO��W�������\L|Pxٮ.a�| Q��u6 ��#�c?�cb�LN+|�:'�˫0jpe�M�E��>�s�䭆�q��	��q�lҠG[���o�Ev��_ 14݁�����X�GƷ��1����������SMBd�A%A���[׈�����'<JeA�v�k\�U��"T�7%��e�%��H�l)��2�j1~��ڼ�g� �����I����޾����4�����Z� b��,紻�'Ze�~�p:0�	�B��Q%���pa�����G�"�A'�~��x6�2��M��(�C�Y���g]}�c�3o��rɵg�8�� x����J8�235>��c�i�|i�.3]�!�:yLy��9�zG�o��R�\�D,��Ӈ���;Tз���<F*7����l���^��J�X��)d����N.X?�y�%��S�h?��)u���u-Y~1"�B����?�3eLES9�A5M���_r$0� 54�o��ḛx �oH�ǌ����ݴ���$mn�$�tB��[�Eb|�v�	���
������ ꋕ�0���7��-<��Z��y��9,RY�v�Fq�������Nr�$E�������'����PH��l�óO���OZ@5f��FbG����u}���8c�W�������|:�� �f����+���K�Th����k��GM�R� J5����Ġ��'��.A^������,iY$^���g�=	^!iB֨Y~�	A��J�8z
�4Nv?�����*�1��WZ��,�xEv'��j��/Iyױ���-�[n�3'���kݚj]�-l����4�cTJNM�f��Q�JG�`ڢ��-��n�R�D�XN�����7�>��!�"��s͚��2O����S�0{)��7E,W��#�t�L�*�6��� ���t|i=��@GrP�a=�X�������O�����IҀ��Z�UbhR6����a�M9���Rm�w��ƭBaw�5����r�}9��ӕ��*+Z��F�N�$�`Da��g�=�*\4.�N��F�ƶ�Ax9n�v����c���<,��IĀK}�uG�6���4[�q6�r�59�Mn��nl�/s�B��m(t(���;�!k[x�\��ݦO�N͆�͸��)��>B�����{�(va�#�C�0�֗���D 9�'��b2W:Mh�D׎���c�X;l�c�hg��ouVZ���C�F'ʙ�8�ɨ��)��P�}��ۗ�ܠe�wx9݅�����l]��t��w}�n�R�Y/���U��"�e-��y�R��*�Blgg�f>��*.f���0݈�(���*�ݻ�3�~HGLb�����ȱ�@>���x@���~)�e�"�P�LEc&�,�#v@�H$�p��S��xql�ۢ��Ձ�/���V�*��<Z8������_���r|��C�@�H�Z��qXB�>�(���ߒ�\�@���,����t��D��#C�=�����ῡ5�t��E��q� �>��d �e��ذO���^� ��yY����ľ
�j�{d=CRꎜq�XL���/@��S��_#��.�����h�x�7��[z��rS�k�\H ����J�إ��2;��M����|j��8�����-�/���rT�Eh�ԣ`���Q�����|k���#6mH7�.k kQby�/f�CNt|����gXA,��j�P�� H����H�'����)���n��&��9��!���d�KOu�6�ĵmu��n��`�Ӱ�k�!�s������=��l��� gA���*��Hlvm��v���Q�@�k}?�[F�/��"���p��z�3"�Y䘌��з&JL��@�I'Rc��T�}�����/t����m�H2�rU�������䀹>�	z��0��֛��NXSPgw��?`	I�j��;>!���d��A���Rҷo`%g��a��B3�gFV�{3��>4���OD_t�8�^��G3����3�	��D�1g'�T��bxU\H���Q�� >F-ĮnS���` o@/ʸ)o���O7��3�ه���?t�T��������р����<�\��0,�&2�$��i)��@�ҽA�η�;�E�̩��b	 �����NX
"('�/�'h�V�yn����%q�T�r�Q��E3D�ip��P��S4�B�T|�J�W����������D��q�$�ޮ.��yF��Բ�n�zc}�C�U�G_�<�S-���hx��L?�#�J�rT�������6,ׅ���t�74���`c�VO�zC?<y2����˓��.גX�C� ���W$�u�����B�[�������`�E�B���&�	.;��
Z�z"p�O�cذ���<��շH��/`>I�����l��ڡ��̦���g�d��$�&�ռ[��Kڔ���~�*�(��o��pE)0�j�T�u�����xL  ��B.s�EEz6�P��?&��KA�����c�I��~�B��H��H�Kò0f��Rz��x}	�h߫k��@B�v`��c5+(U�����(d�y��SqL��Nm��.QT��qV �GdN���y�N@��,�6�������y�0����OB+Ya�@��p�{#ZOlX��__9�􀎼���[��5��b�&J��r���l-\S�����Xd2�u�0�].�\���8g�9Ma���pN̚QD�U�n�}s�:?j�?k��H���\�9��ݸ����Q����N�Ȫ=]��\�q���U����!n/��A����<C�'���ӛz�]_���˅���!O!?_����8>�u��f���]6��̔�W�.�$�F9�m���i��|V�~0͍��Q�"Ɓ"( d��,�u\6��X�~'ؗ�#�?M&]%6ڐ��V�9���A�4�P��`4���Myb�/��B+�:���TSh0�g9g;�<Mu3�Б��T�7�:�(�fB�Lw*��3�G#�!$��w����Մv�����4��g#�Z����Pˑ��]ER��l�A����W��ł<�=�6C��/���U_T�R��Ò�܌,�iA��䈄���8o��I���u$����
�w>�����O/0W+*�E(�l�BG�I61UQQ�>[wUCn�eNJ�&���^I��g\F�X����������mu�?��Р���0��:W���K�
>��z����5���(��eZ����Eհ7Ƀ�'w�(]��x=^�0��P��So`^�Z��<�D�f<������b����[�lq
�]W��2����̍C��z�UV���G�K�J	��Hs9(��y+c��*M����/�p���	,���Jr_���c�wy�U=2��4�U�"�b�y�q*�?�E1$�|Y�pV�QF�R���9T|
L^��l>l�?R��O���E��M:8����- ��OY;�-�H�,׽a���_�����J�K�C�&T��$��Q�r����w]m3���)=,��B聒��3
�N�A�� �.�jdg�0�f�6.��:�S�	
YZ��z��LC(Z5qz%�1�@��K���*l�����������Z��'f=� t�"U���pT��ծ�k��c�(CŘ��%�°ʿ�=���%2M?V�;��$�T�ܢS����pA����]�J"�◱��2�ɋu�0B��Ib^4k�����p�� �Zz}�t��P~u���̷o�9m2��q�!��>�I�W��4�����������+H-t�!�_�W�C
�I����{SM�}LB~QB=<q�;����F�bٍ�3�h�� 3w��և��Ϧ`�����?Џ=�Si���QD7����>)�mx��jq�Z��@(����]��c�z�i�re�Ċʪ�쪧�_�6�7BU��%�\�ڟM|�qP3����"Rĺ0l�@A���@.$xSX��Щ�����fk�>�6=\��ojUR�09JQ�@Y�v����F4._1��j�}��<Ԙ<ɆW��5H�	c0�_�)�AO��Z����9ڃ�Z�ؔ�Z����[<�Xl2z_����K���}�yV�1��ʾ)���X�����+��dׯ�ý.X#�,���%m5c�+��y��4O7��ގԓ��v[��l��UH����������ƪ��O�!�[Zjl������X�X��G��4�����^(���kM�ͱb��T�����/xG���R��\��Yx��QB�mo�뤭�� ����fy�k�b
���*,�H"-����WŐ#k:�P�q���0/��A�韎�Z'�ܳ�O���2P�u�q��}���b������4��=�0�Dbo.8p#��]��"��>)נ0���q�k�q��^�J)�����S
N�ϪY���!�TU��?28���������
Yi�d�<m�ab�4--Zd�'��)��|�o�'߼��K��~��4qh��/�ִݳ����'$1E?|G��v��n�B�:׍s;Ѝ@��l-��'CysP�K@��vf)`q�u/}������I���֊��'��ռ���c�CqU�w��TJ�P]���,�������I��Bd��Y省� ����H�Ȑ���^�����Fغ\���h�I��Y�-<������x��dM���|Z�9H�e�*�uA5[�� �y��~m�=��ڋ}n�IC�|�$���]2U�(��k_;�o�ip�q�'��%5�")h���sU�r��JR��s�y�
F�c����Fʤ��Ԃ=�m�B��V����� ��F���sq��J�c���94ޚA��6��5�zV\Ki�ҁW �,����^�txtt���@�Gc�y����	���P��-2��/U9Ra����tY����}W����m����]�F�vw<�خ(�:A2 o<{Ɇm��4�n�3��Bm�_V�������̂WU�������Ng���d{XG�߹������k^F����^(w�s͹��W�甔��tV#�E��<*���y�����hf��(����I���ࢎ\�Y���q�K3�3�_�������R�����!C�|�ƪn�sZݴ��V����9ޭ��o�V�L1������a����?��wD�^2PK�kSxX΢��Fx�������޿!%e���[h,��h��a���Ɯ ]�+��#ɫG�Dڲ0<,��,-���/�%��3���X���"��-��`!�������+�*��~ц��NۍW�4|�ggU��C��T�^��F/����]y䘸�"�"�Z��NDF"'\)}��#�r߮�����,(y~||įS���/]ewE�����L���&���)�n{8�2h�$�ؼJ���<~)��R�YRnq��`V�/�u�HS��wL@z��.�j� 	U Z���ʎ��l|mAϔt*y�*Н����'�3�m\l�e��j1�<mw�T���+=i�6Z��R���mX)Z=J��rgDx��_�35X;�o�t�7�w!�6fQ�&=����}<��G���H�	�B}��� �`&��]w~KUN8��z���k�C����j_���ա��aM��H.�j�f�k�`eyP�6�fx�T�Q��FK
z��V��䉏*�O�v�1�("�<�g�97��,B=�������&��u)) OD&_�X�哇*�k׀�Y�u��1ׁV-Xe]]�6�qž�h��f�;��(���;|y*h ��b�O�ЂQ.P�qc"�^�c���?E� �<��sb�"c�\wn��r���I��B���<>��j�x�'�W���T2_kPkQ�"�|%_m�+=��z���k� �7Tw�}E�Ȇ#	�W�*��t���	6��K=��s����E2��&����Sa}�w7���0��:b>=pmJ�(�P��xK�;��]~,�a5/��9�-oLSZj�L��X�#0EG�D�i�ל�B���,%
u	T����?D�i�N5 ��팙"����赞���B�$ΰx��f����v���kD�{S�˅�>Bb��ˈc�~ẻX(G�Ά����h౭�s���6�&xŜ�����~^�)�<.�*�'��JZ*ܚ'��'�m��\w�C:;��&��J&�N�&�v��r�P����"'���8����;zbH���/S�<��ږ��GK�y=�DV�Uk!}ۺb��Ң�҈�PT��-��/Xx��#�Cp^�P����q�dƎ�ɀ�.J��9 � wH��֍��y\� ��R���m�&h9�����$@���TWЧ���Ϸa�JJ�	��l�0n��7�\������p"������m4���D-�b�	T��#Zw���&�@��!@���j��&�����۷h]D	f}���j)�?v=�s�@���w��M�G��]�%�D/�Tz���Thu̗ǒ��k�l�d=`�9�bI��R��QPl�_Z�vP$\��O3J��2���^�� �߱X<�7��C�Vp��;WK��H�����(��e� cr�[��<�U��������J�-��d}i�wqQM��vؚ�\|�#�,��9QI8�p��V~P�}
�8��^2_k���E��r��α�HG�5r����`�?෶ˑÏt���W#�vf�!*ͱM�)>��duj��b��'�[gL�Bb��G2��z�l�fl�u{���U0�νl�C�3O��®^���4�+< x[�Q���^����?_�̽{�f�n��/K���+d���j���N�ŏ�T:+6~X6�E� �◆k�zԉ��l�#��&��= ���3���=43.}!�$K]h���c9�3+�B�+��S����Y�7�j���"�J��Ou��sE��m Eҗ��y��k^�.B�L�\ȕ�jMc]��H����_UZOk�4�����6x���LuW�E������!��d���Mc�tR*�QNW�䂻2�3c��T9��� ����b�j��,����AT`LmJ�$`�����
�
�����b�m�v��;��j8gz��!=0&݌���bk�I�U���B,���^HsJ�����Z���)`�Q����H����2�4��d����N}����SC-;@�	��b�8��*ɭ
o'ڶ#�(Z��aO�$�T;}�C������?�)��S�;`71�tٷ����������D�#
/t�3��KDc�7��'PY���O瓚��u�96�[���6<����SB�]�^��܋Gf�Z 08,F�1[�>N��R-�UE̮#h���%r��VQ�ࢴ����uS��Z�ǳO�Q��a�K��~����6�c1a�@׀p{B|��q�?�Y=�7W�g�T[d�;:_l�xv�'�ޗ�?A����Ā+�$bm�J
�y�̄H�� ��*]�	�æ�C��[|��}��0�r|n�$���)7��4��`텟)@Qo`Tʃܜ�_SL�h G�,oy�3���Ctv����n�\�~��]��#�V�p�9$P*������k�>��4H �I6�{�8��-�2�Q��� 6�ȓ��a����i�<�+M�j-h�=Om騥�i|��/�
����p'eMZ�Im�Trd����VI�aNO<��8�7���.0�Lmi��5��
���E+��O5pvf&��p;[�<��B'2Z��7��� ���E�Tw�WWC��?	����.�	�UPw��M���y�B$�/���=pj��j]�*זuHؑ^��>yA�MYtw)���zV�"���/Bea��=�jύS��N��,*^�,�Z2��S��R��������y��[��Gs<���ɰ�b��o1���s�b�Htj5Cwvs�Su�l*y<��9�~���]�U��ċ_��Yc=����,���v5WG��s	Y�(/3��(ܢ����_3:�,Ƌ�o�`pW���˓|>Dg
���tjMM[fbv��)��F�8��Z��{es��X�z�d��%���0��4/_WY��x�� ��m�n�E:��x�/����oW��g�������
w����{iZz��l�r)�3Zp�/��@����>�~���۝&<���$F�U3��}V6G�É���fo}�W�i��)
Z���4E�Yifv��ѕ+F�Z
�����r�_P�8m�L��R�w������snA�[֝Y2�m�Xi'JyY�q��YVsMa�=�-4�AZu�B}i@���W�!<2�y?+�{�!�����X��՗V���/��>��IL%w�q礼+����0j��gb�a�W��@���U���39 � <*�}���7g}���<uij��$W�2���m'$��A���8�L1�E �[ F��k�.�͕��R��1��9�o"�t^x���j���T)�R���7}�l��Ϊ�e� =���JK�XL.%��[vuH��Ԉ]�����䃑�-����v�љ� �cħÚg-��ǛE���ɭfD�(��T�����Ǵ�1�K�cB渪�,R�f���2�Ml(���;�(��]�h�Q ��%��RJ�Մ���xD�A3�/��FIe�C�	���P�x
gv�E`Y�E�%���X�z�c�D��t�#������&zN�ZP�:�fP>�X/%nS��t���y�|��Q�+�%Ɉ���_�K*sf�]�(�,5>k�3�Vݚ�f5�X3�����H��sg��Q��e_�g�@�潚ɼ�A�j�`�!CNYh@��� c��mg�nS��_�Ñz�}-I=3q�0e0�.j�����K��aV�Y�ۑ��Ua���k"Wr�Q�I��\�@��� �sH��-�I���R�
��۰T0�n�Z��������ּk<I=���H*�s��0p�I�KZ5���ʻ�^]�d=�Zp4f5���������ǌD��S�zS&cp�^!=j�[i�ٮ},�+�)��zlHd ��^�1�~��|����X!"�k�6�C��/���A�cc��D���A��%�/4�i'�yi�a�;�b���<ڃ��x/:Gڮ(�ATMSp�A��b&�e���$/	A�/�(M�wo7����Ji���2X�\�q��Չ������+Lzq7�'�Hd}�FǺ+����w��l�� ��Ǆ��k�&��ٿ|(�����5�8ڗ�9ң�;y��'@#�U�>�y�����8�c�����~�-��#����F����P�(���P|r�D�Ś�8���#\��Z��O�S���"��wRM�)G���8�tA�{_bQ�w���"���E�Y�&�ti$��I@���!���
���7M�N���W�� >?. ������
Ƌ���:�ZE���r�r�ow��hA���Σp�Wh
�D��d����K��`*�P).��p;$��FjF�F�|�r�i3<fŃR��xF�G�p!�!��f���9Uz�GY��ל�x	���R���ė�,���V;򄹅��zW��TB_X*��r �=p�Ka�dܽ��m�t��P_dL�KyDʦ1������(��W�c[h��|O����~�Q��y!e��g(�Hy��G��18uJ���g5t/_2�j��U2$4�S�cJK�5@T;!�� ��~l���&��3X�	ׄ��S��:01B��p�j��)��=K�Z��F�r�1K���d3Qܮ�gn���-��:���U�@K�t'*x��3*�G�0&�y�0�^=]����'�;��z�PHC�����R.k7��);M�rj���2�� �@�6TeZp�pу���(���!@��㛰 P��q���
��ۺ�afq�ʼC�`����>z�
T�m(��5�s�l��f��%S�)Z�)R>5coå�8t��b����p��Q誂���p�/Z�ʹ��&ԝ�ĺ�_�C�ƈS{��0�(	��B�<>Fg(�&�b�w�3��d[4�Ie�<gT/�z_!�G�&�b��/v��A������Ak�� �Xv�����J����� �x��p�j�>lcO�t:đ��Ô�;���u�U%�%u�Yέy�'Z�>�	N�};+F�Q���Y"'��N�nj�����>A�2��I�)|�HNA��h#�����0D���B��R���{�3h��K�Vj��1��^����)S��N���J���G\�t$W�u�l>���;y���P���I�F0�7toɉZ"%�W1A��Og��g����A���_�PM��/��=t/�W�L$�z�#�Tt6��]߉ nQ�2���MODe��%�}�y6�a={���F�*n�ra*�����`s��-�P{�z�q\6Î2�����+Gi�YhОe���`���������R7��E8��ԈI��w9�x���,ƹ����ؐdzk{�/L����F.�c����&�F(� �'�G��(�S�W�"��n�W7��r���=L���ۘdũ�j\v.�oC�h�{�Tc^*�R�b�$��
�T�p��0��m����`���?GÒ�^�������_.�
�;6a\B����C���?�VY[��^4H�E��g��%������ͩD�g���Tup��w޲D�����jQsq<��Ī�L]&6�����X�v�d?	Lo����2�,�.�����2<jW5���l7��[}�*#�BAfr8�H�8G�6Ea�fv��J<h3�ָJ��]�,�YBT1/��A��mF2��Ύ�
�֜���ݥ�����L�}����/����$L�Үl�䟥B�|���SGiM��ů��%��y5�{]�V(~a�n=i�H��k}C>�e�$���;#:z�
ѱ�{1�p�Y�9a\��x�	�6e+}� 9!�UEW�h��#%�A���4�Rl;B�1�f�_��s*�%c����)s��9,6!�1L�6E�L���ʕ�r��6T�����s�E�j^�˴o���&�:�� .�3N%���W\ N�;*\+Z��(_n�5��_�P��A�b{W��
�7���<̹ՠ������F�gŲk0�%���z~t��!�\~v��ܯ��7p%4k��K�|r^�)�َ3�u~���߱l�7LB�9���^�((� �j�A�v�����Vη���F�΄��n����ה��#�ס ��������1ѩ�Dg���^��-�J��K-q
!kH-.�X� ԕ�n� \z�s�:qlɞ�WN�&1y�b���n�2R�|�Hd�+N#N�T�/�9���Mg��2��R���ǒ�SIfїy����_-��]X�	��\��AsI`QQDTp͛�q�L���b�p��·�@�d���>��ȸ�:�}�Έ'��hh�Tn��c�tT�ע՗Q�(i��*7~��ه�1_����(2��i�	��
�AN٥�o�	�Ê�f�������J����|
}�A��[���øΣ��+��:�`ƕjgR����V^��"R��h`N�Fp=n�ٴ�M�.��_�T��˵�<��ȰJ�e��o�d��X��	~x ���2�p�'8ՠ�)��G�fP���*r0J	�����յT�5�ގU���w���1���`�J�"�I����8k����{�ﶤ"���Ԑ����������S���mOœLyNa����W�a���$��jn�g�逊���@�W�iT	���ӽP��<�H�=�s����%'K皋����ڭ^�쩕p�U�BQ/x_2�\�#��s���+37��i�G0�n��������5�4��)�#�����Qx�VI�|i6���rÚt�`�qzrs@LC~�
��pQK1����/�@�⯽�|�>�8�U-�h\.�H�'�j��UK�꒮�!�[���b����}��'~M�i�+8�1g��1��e�-����Y����ہq�3�cn,k0�H!��__"23�cXYc]�xM���r��W����M}n T<�$X�ō�U��bp఺ƢMk	Ln�����S�.?�0�D��a�D'�b1���)~����� �D�l3��Z��M����D�=
\N�>,��ǭ�Ul)�U�`��W�~.w0qϢ���)Q�W��c���ZK�rO�[�b�Y��[��T䋀�Ǔ�!b��wP�EgZU2It><KI��o}[HE\0�Eʖ��{d<d 73ے����� �Ƣ�!Ͻ�ĉ�oL����c���8�[,���%����5T��k�DX(¾}E��M�d �a����&��2�y+ӣ��������o�_��L����Jχ^�R�}����2��E�j䩬m(��n�SJ���eK<M�h�D2
QC5b��:
Y�����l���אH�E�6Y�${�
P��oc����tc�7&[�Ɩ�I��K�|=8���ܿ�7�f9�C�D��k8D0�J��py���Si� <q�{0�6k��ܞC�T�  ��{|F���) G�Ԇ����v�G�7n��9��Z�+�J¬A����B��̀SW	`G9�fj������͝K&��v�: ���5=��\!0nR�j�R#�ѡyJ�aU~t����=�М�1�
]��t�K��d߹�X��5]�a g����VK�od&�e��paj���s�m�K!�ip)VѮ�3�5�g� ��>cJ�����c�� ���u��9e��%���7dþ߹pڻsum�9{��^�y�:�w�٪�)�ƺў��OC�nX�v�&��s�N�c��2:l�=��KB_��hfLˮ#"�B�����a�<*?Rn/G|~h-V�=��F�@�2S��r�qS����p���?��l�{�Ow�G�=�K��r��^�y0�`�qU�6M�0���F���z
3����8c}�Ba�T�ト񞁧���`?��a��:�-��E.�6��ʅ���[U�CX(
��p��?���F࿍c�Ϊ�}GĪ=�%�:N��
T�I.K�P8��i�a������/h��\p!̈,��,�^�"�VNp�@lx�m<L�
�Z�A��MC��@>�t~�L�Fn�=��P�iD'2_��2���1���e Ư�J��7�'�$����z�wd?�^�0���s�*�h��L�V7e#�Q�!xx��4�?rt�F��J�K[��fݖ�]a�f�D�}6��x�%� K0B0gJ'u�(U��xj��LP���x	�#��Ͱ��V�[�j nO�"�SV�]��oCo�U�uT-*l��0�Ί����i���nШ��O��RYL�.2�p�(�0��n.y������&i�Y5���I��l":�����k�IO����,�A ��s�X����0OZϑ��v5H5\O2�
�|�P�儸��n��A��N�"��j��O�.}Q�(F��0'h���3c/]�����C�s���k >E7�w
�&�0�����1��І��h0c��	�+�H��K�l�i�5��S�7��h��Rۣ�#��;RHB��#L�������5�FzO.��,��%g^��=wN*�;jᏰ�ѥ%�)\� U��e��3%ru�nS��������X,S"��/!�E&gL��)|���z�;�R�=��V#��k�u�	kC����C�ˠ#˙N4b<� ��Y�	�!}�L�CF��1�����U��?�1��ǌ�I;>k%||��|���!-e�״�K�Z�F�\œ�����a�8�8�𡊹���c�`$��O~�^K�fά�I�ni��I+��,�`)�\V�b�9��FW��A}�V�%�����ى��࢓��8؝�h�@�����݉����Q���qt�ڶ��q{*�����i�Q��������;R�|ô�?�C=����oF+�ҿ(5��-CtY/��3�I�aS$��l%��/ڣ�KWۼ������8:kj�V�^�#r��\�
��U�7�aG�E�D����ep�K��>w�T:�C��4���]kXQ���7ϗ�W﮳>A鵛�=�f��D;hV����K$�xx$���	[`if'���-�%T�
�,�>�Av�kĬ������ҹo��r��nL}�T�|�}�}��wzը��)ؖ!u3h��Z��!�n0g�ݺ|�^�g�r�_k�{!FLf�͍t�4|�H��z�c�U�}v�p�Sue�̚>�y�l �zM����x���6/^��ZZ�<�:V'@���1�T"�D�9Zh��MS.<+�֮�d��p�/���fh[x�� �t�;��0�޻Q���B<�i��o0���|���f��ؙ��M$�	8�����w�(ʥt� �iC2@���G7򟸵�����zy;^�RӀ��Į+$U��&��ƶj����nC�w�M�0*���T<�
��)� Ș~�p�� ����"P������A�5%58 ��E}��֥ ��/��0�Z<p(]������`?Q���5���;��}��2���1U�� ��b�~�?O*��Dמl������H�������JL�*&X{��1�Tp��ۋ�$�������<�>k��89L*JK�c{&��]�]wVd�K�,i _���N�v!N����B�|�&�d��(� [~�ކ�n�n��Đ�RY�c
ؑ���G}&Բ��/ј��#юQ1���n��zy��m!8߂Bj[| �cv	���Pwы��l-�M�H����Zڅ��wHT��u�Ԙ�$���fݑ�Q�Y�~�����l}_�,���,��@��ä�W49i�0x��"[�R=~�������BQy�����eG�6<ޜ�Z/�s�"�,+���rp�qorˬVn��H�<G�!}��X@�T�Ǵ?�q�c@�k_�DXXJ�����J��A�A�V�p�yE
��d��]��k��Q���ƴ�.�%{�����A�I�S�u�[�_���x�n������D�{��MO�v�:w��֜Z�\�j��2E�@@����H؊]�O\\h
ܮށ]�v�iv����׹�~H�}rtC�g�[㇂a}U�Y�˷yg�w7�ɆG>�<	�n�;�ld�v��@�I�~�u�kR��&>sU-n�T��h��ɡ�C�+p�d�#�]rށ���X\�(�6���T?h��,�!5���ʷǡj!#�PDo�5q�^���Ba��*����IsmVv6���9O�+�<Cyc!!AHDI��e�!5@2�{�ձy��<�-�h���*o933,�CWB8TC���&	;���n"]"��#Y������b>�����2�l���*n�ޭ^M����W=n��֒e�'%c[�"i��<���5�k����H�(F��e�w
:~y�Z�=���n�*PB���
G�9����W��̭�ni5'��I;��]����ܾ��K���# zù�&E��}���O0�ڥ�S��������� �|��h3�ۨF���E�`�!9Q��D\�������G��z�%����P �S�g�3�y�)�tN,M���L���!6 ��l�c��7�7%�󤋍sT�pH5J�-�.@2&�����k�\�S��l�2�E��|`��b�yL��"���(�tc)��f�%��;�4bw�ky!S'�	�_p�.���X#W<kdlr�pc�Ңqw��%nF\��g4޵&�R��t�d�X����6o����!z�
��������|Lp���� D?��q�LAwݢ<�����gE�i#�C����{���D�p�A��'�74C跻�p�*��R�4��2^:�g(�Oh��(vw��O��o���2/=�'9}%���mnD|�>:�Z?��@��H��7�K�#�Ţ=~��7��~Ga��:�6!�ǰÁA�ٴ'W�*���Zƴ!]*P��yD1���_ K���(�A1�^�]�����F�ø��X�v��Ϛc��<��?�j�&�A7kV0 �(��uӠ�Sqƺh4o>:�k�����8mT>^Fٟ5������o�G!Œ�ՉK�aIC�á�	!�����K�0�_�=��r;�~`���*Y���R��Y7ΛG9�F�CQ���a*g�x1�U�/�V�J��$� �����:���:1�K�$��ى�)8��
�SC���R�<�e����5<�l���.1 �!x(�![#�"3ym��H���MH6;]��D�C�aE/�澌�~��&�=3�r}���3U��s�t^w}���n�޷M4�W�����ܒ2��p��Qݧs�Y+�b��ϱ!�����8_��ٌ�ҁ�����2\ҳW����SH���� ���c*�����W�J�^�	���aZ:&��}ϑt��F��E�Q<U�٤�� 	�cTg��6�|�w���-�~��e)����/�aS@#���>��x�Ӹ�YW��-�r�����؇9�� E;��,��
s�Yd|P�4+�,��L���[b]���C�-���<�\�;������c�ۖ(@O�#D��[xU�p/Z�5�H�a�L�sĜ����������JO�(d�kF٤���C�;r��V� ����
�]��
)4w库�vR�RsU?.��[oĥO�������E���o��輓	Q�.�W��A��-���h�y�CJ����~�;_krF��\��YwkeP$�:�͂�q��W9����2�Nk�(3@7����C�������B��X�#�4��������#I��N� �E�Jxh��H1p��q3��H5�oy0d��F�	c���=�/mZ�,�ڵ�D��ˇ����aH;��s��%�iB�p�m_;g��TG��@'��tw3���鲵�Z�"�����ս�d�2��O{P-�� 
2{|j��6ވW՚X|@x�pU9O�:m;d�}�3�ih�_�q����c�i�)���,rl�s�-��%�����9���?���RəR���ܗU��>�Ϭc�LC��M�c�j����G��Y���١��=�B���䉉����ԯM�k�h^�:,C8�v`�U�&�t̛����޹V(ʬ�OK�2ү)2�n��B8lL�f}��M����K��9佝T��?f����/�.�؎��?!�: P���ff�q�7���a��+�2t�m	�_9\�CN����[m���5�J�0���Ӊ�l��R/�?᮳��Ā(�'lC-*�3���{YãP�/ڧes�1�I��a�T�$N��M���2<"Z�9~�9�Փ�����/��+4��������1�%��	����]!����r�쓼�o�T6�NH�MR��9xN�!�&���`�M�U&��?��+�Q�Le_�t�<�i�Qb�^���+�� ��T��X�77-홆M�q���� �8k'�aH�7�Qnħ�r�O�2p�:g�o"˧��f�H�ߦN#RV���_|
|z��?�$B��7��~�_\�q��Bil<��P~�8��2#)C�)���Y��..����Ȋ��'��ܚ�{���ͧ�erS۩�n������po�\�{W��徢N�~���KJim��%���Adp�*i��Vn�R'	NK�[����ҭ=T?�2�^�Ī�Ѧ^�0
F\rCtm��X�����(�7C��|VE�������ʹ���N�}�_Bc8�F�7GR=N�ãf�U|��lj������p)�S��k��{�,�[�:K�%�$.5�\�!��%�H�*H�+M��1 �m;�������>'��kJ��8��6�\]�����:{� �K����q�bE1�k	�3��[l��v��
}��PDYܓ�~���<�H�p��f���)��e�z�a�����#̎x���ڒJݙ����L������뤦����&��[���hT콅l
���r	�*-Ӂk¥�Jh������h�`��URu�fp�$M�����Q��i�� < �K�e�v����gJ ?V�f���h�lW����Q��g�����
�#}w	��s!�k9^f������\]��FQʛ����ͅ$�	�]�9BIt|'9�Fp�:GRg�V&��E�� a�ʟ��;ڴ"3��S�F:�`�� D�hZ���P�%��)��5��
<=ZK78��{�=H�С2�}m7�M-�
>��)9D�N���S0�H�W�"�ֽC>Ljxb%y߱k	� ��>�+�u��F��o�o�2�����.�����Z��ע.į�90��?�(&JK�s��=�p>�~��F��-�Z�V8:*R˞H����XN�b��R�#�����T �a���
BPЦ����-�(��'�P�G)Y�U��&��� �by�1W���n���Ԛ֚_�W��Qu2����L�i]��E �M�2�Vwr��]{Y�q �O1�Z,�3�Z*
��q/HER*�ȍɀz�k�n�]>��9�K�G�����K[_����.r���?	�{-������j�-�N�<�^7���O���	u�0��X�ItKL�~���r��Ҫظ(M��fj)�0�����k�����f_�hvT((�8ohOFLQ���~l�qK��<woDߜ{�"No�xn�hKH�Ҿ �&�|*.�>h���<�L�|}k�bĨ����M!LN�H�1bGw]��䱊�^�B7u���b`ON=ȹZC�Ϋ��\a��=\��ړ�o��6���;>�ȏ;�,�u�N���o��v�a���ߘ�*'A�OCJ�����'mp-���7G����/�w����LR���̸q󧮉��-v�bMQ#�t1�����Y�^$=�����3�dSg�����`�&h0l�u�Sq�ca���	s;,�ռޜ37'�5؍�XWF�q�:E��G8�1�E��s�Y���З��(~������>�)k�ڄN���Z���b~�AlP�gyZz9����S{_��l[��-y��9^�#�	�N�V�e�4a2��޾H�fZ�K��=N%��Qb>��(�Xo�k��c�@&1�gQ!B�|z� k��6K��|v4�|��� �~C<��]ȅ�&f�n���h�_��Yd�/[Ɉ_�b��	�fc�~\zF��e2h����`K�+�-�ĤX���N�5�ګ+�j�e�����O�9��!<��P�!6r�Й�Ƀ����uv�[�#��d6a@��0l�A���b
L�/7��O������*�!3�3�vl[��i���3�	߳���L���17՝۾h��l��S[C�U{����7�;T����l��PF {�M�L��� 6zNѶ�hy76~��k+�nYق@f�J�''�=�v2�s̪F�(ִo�{�3�p3��7�@����X���,ҹ��mP��1?~5�ɏ�ˢ�b5t#`n��6-x?7D�ut�5"[��<axĖ�A�6l:qZ{�����SDL������cU�  ��x�W�q<u�[K�7l��8��]��k.�
~9�a�n�:V �q�}�#����`
�bo!K�!�/� ��d2w��ᠳ�d�u������7��6m�Z)�RnzU.�3,2�f��lKݰ���Є���"e�;+F��n8�E��k�,v�̉��(I��p�ꡅ�K�,�E���OY��Q�����8w3��o��V����㘒���.l��>!������<��B����%A�@dB,�����Q���
/T��H@œ�+#�QL3A���C��M����yU>iz��햝FF�|?�?��N!=c�6rl,z�)2���,���gE���:)�!꒗[���ĥ�9�J����ms�vT]���$o��K�I��°09����p�@�]�Nb,��r񶜉�!k�r-@��.7ë_υW�&�F����מ�۔Y]��f�W��r	|[�Ԁj��V�����͗����~҃�Rӻ��ǟ��8P/D���(�U��s�X�+���~�g�	챫_�V�5n����T[H��1�O}É@5��[xTM�l�Cד#9���>$��c�$ U��TV
y�u��e�⿪�yQ/��Ci�J2�X�jU������Jq��~0�����9��n��Vz��I��nC�զЖ=�׎"���#��V�OH�Uwd^��̯\���Z~QM�Nu!�C�ST��3e �v���o��x���.�?��8W0n���iC�����0�����YȻ�b��� �AF�d��I�:�O��o�,������L�d\�(�_��� �:���PS
2͗Nu�du�Lco�+�����T��|��u[6��Ϲ������!f��k#�1W�P��I�m"D��{�����+pǇ�Y�DQ�+���1���~�MZ��/N����o��C�����>��۰C���}��Џ��78dt2������<�~ڰ{�%��
�\�KS��l,T̩�&WE+��i2k�b���>>��g��*}�P�|
^R���ů�;�!s�����9�OL�[l$�o3�oe@�kݛ
���M,����r��9ZYُm���Kt���C��;�u1��+�偖ɏ�=�o�9�š9I��5�eG#$��.Č#>Xo�J4��I�T�%.�A9<"�f}�|`v������f�7�J�/���\��N�'���9�����vմ}��?�+"�����}w]��%3�1h6����d앐�`+��i�M��K���V�Jc��@	j�:�PF����W5#Y�=c�Y#5d�y/[�U@��7��Ӏ��`�����\�`6?`��}�����f.���A6�QA%=�eed�R8�#�_w�Ҩ"����Pdݑ~�������o�Hyq�y�5��۴��׉4���]o��-c6g�O��K΃"g�s���R<Ѯ�t��;/н��_���~�Jb����b�B�4=^�ɥn�-��H��K�c����_����Qr��a�<��u���!�h)Dp$���dȖ�m>AP��D�
N���-����99�LN��c�OL�2m^�s3μ*1k�E!{Pn����K4w[]q_e��������^�V�c��6��-1(��`��Tl�W���}����MD�^��7�p���,Ӫ)���1'"���뎱|Y�
f詍��/�,�GA�f�����j�O0�
�y�ɨ�ũk�$eZ�������\:Ӡ�kZ���0��-�7)~o�#*�׶\�q��T���AR'H��A���NQ�^�N��Ǐ�y�7�����;�����e�a{�A�ğ���Þ�r��kU�𾲲��`�q�$�5Ť�$;?՗�H�S
��.�O/�T��܁C��9����y�����g�:����9y1�T~��g$��^��{#��l5� ����,�^r	i�Q����"� &���

���ow�a]3h��XR�5*=F�Hi�n��U�څF��V���C�'���I��S�����N7�9������j���|���
>H�6��~�ǜ���nf�jv�s�#1�=(,�Fe�g��mѽS���n�����N�3^FD��;�]!���}�������"�G+�(���8s�."�*�&h�d��zF#ưxy�+8Q��6�8wKX�"��7 Ƿ��×N%#6-��Cq�!b�E�RN�-�����_N#�H�rZu��)�N�����u�n=@ٟ�[�G�<������Z�G�i����4)?>�5N��M�Ic�]�v���맟R��
6ɮ_�����O���
���j��S�߮�܁N#���6��'�:Y7�cs��h÷S�Ft� ���<J� N^)��N�i<�Iy���Te�{��i���{���̯Զ�6c oc ]�����v'�xQ�ٍ!c�Vּɱ<������13�u���u����,�C&�ٓ k������x}������� TU��F�6s��|��؇�K���q� �-Fy������f�|�����ĵ�!�;��E���=Ub)@!���r��'���R�^�m�j�\u��bo֢8B}6��9��=2F&����,�Te��n���7�x��	z���u�е&���	��PqdIVN6�2��aU���7�J_�0�B}��2�'�}�g��V�vi8������Go����͸�A���v G�2��'���c�酇L�v=)�kh��-8���S�wף�&d�Sڇ�e0���̲*���mjhM�y�]��E^T4�0'��Ga��=�x���?�Z���io�+{7�ʋa�Q.�Q��i!���c��b�$^�7���6�����X��6k:�Y����S��K1�-�+�M7�V�0��e��*W�QΏ&w�V��4���'H�8����5g�LI����IV��O%\y��w�~juO���4J8�'�i���ʂXy���Q?�o�Q�,��=/ۯ X��	i�hp��	H Y���D�9�.�O3� {�o�K�s��zZVv �]+M��P�R1�/ĎQA�d*��e����c|�b��=�D�H'�K����6P�3�0K���}]�&�`WCZw�|D(��/�Ay��ג(nϊG�ǟ�M�dP=��Ky���6qjn<:]��Nr�ދ8A��B��"�.�Db�E�=Ň��w��%���t�r���lb�O�Ͼ�0���R%uR·�@��`��O��8|�S*�L�.��"R7'	��ʻ��\q�������sM �4��:%�"kʙ��3�v,!�$�շR�fQ�AA�n��I����:'��3q����@��q+|/��>�2��g��o� ��E�Ka*f/Ex7�H�^��&�a9i�����2h�IȎ��l��k�GZ��B����}��~� ,�[਀+�z��(�B�H�C�RV^Vkk�u�G�˱����ק`edʰ����?�z��E�aH������vI=�Ok���� 7����
����M�H��;-�!z_1Xd$��/4%n��4��
h���ϵ���3Y�r[I�Lร���R��O�j��YL�!���q�w����8��
�� N��ݜ�f
a��Deg\xJ�a���$���}Z:�vx:��ed^w�o`��K\�g�|Y�3���+(��������V@��F߂ `j=�I-9nc!x�Pm.f�l���aƨ����(�8���)��M	��v2'�Ap���?D���?@���ȭw�J���8#p �aJV�Q�񇻍��Rgx%�{�
��;2��æH�M�Zq�iȬ�Z0��фr�0���w����D�%�/�^�9˩G�ѷR<,,\Nh��
�\트��8��L�2/�Fs>zd��|��2~���G�x�l�3:�dyIr�`ښ�II5��g��f|YU����q#�ߚ8?����!3��+0|3��C#�����d�q}=x?�@�n���M��t8/��&����2��"Gb3wS�.�9P�����#4���\�IZz!��7��i�/����|���Nz#��p���r���1�y:�.<�r���qu���m�v^.� �rԻ�N�3��n���U�a)��$cf�+���0m��!O)u��~b��B9t�k������X�S�N6}Pv�0cu�p�4���:+�M���!�PZ����K���f�I��*a�d�~��,��D�I�{=�Pf��Z�֙ο˘^!Q�7����Ӊ+���'<gy�6�v<F�>ivqL��M"0}G��Z�,�����W��%����`�w��^��
R�҂}`#�vϚ!����`{�$1�$U-yb�R2���T<S�J���פ�@o2���eR
�|��rw��T��;[�*t�ח���F�n���{ϴ{��ݔ�0���KM�/�\RH���dv?���vcY�m��:���/^�O���]N-��ժ10���MoSt���خ�k������$�`�^�`��Ҁ�QA(��(K؆����!Z�[R5�7�Z�r����[;���^M�������H�YL��C�XJ�3Cs8"R�a���`?�Fl�H���ԅ#N���\Y�l�������]�0h��:�x��jS�[+�)gd|�[~*u~H��& �x����|���OҫL4�p0�C�q�F�h�<Z�S��˖_f����d�v�x��=O��%=yuQ�0������<���?;�2"�9���Źds2��P��F��A�zPe�#N��[�v�����%F�z¸���I��9��_���� �,�� (�� ^� ѯ����O�����k�m=F��X�����Q�8�-����nV��:�@��<#�"�z�IQ�tR��DK��!�)% �����'���,�����6�*up�y]vF��̟V��>�������7��u����ZQ��	�0�U�(f�"�q��)H%m�j���M3p��h��9�k�0�E��źiu���+�*�eq�_z��V�LH��W{��eVm�����j�+7�V��~��#O��i�S�k�R�X�R_2��^w��3(�G��a��x�4՝��#br��}-�ٓk���Q��Z%�<�˦�1���A,ۛ�z����������;7��)D��ԛfh���=��I_��cyD�}���t���tI��4��+�t��9�Q��� P�S����c�}V�l	�~h,���7v�M��d~M%,p[s��n4��?�P��3s��k���b,��Z�q�Se��;���d�E�ِ>�cR7b����)6���\��l�egQ4�����rPc��#wHmPB{t�G\���_`
�z����l]��E�, ��}��ڻ���lS�nec$�5��Y�m����`mzX�8�;�8`�m8��7k��*xL�Ʒp2��gy��"��_�bN���7+��=J3�����6�)`}W�{<��7��\� @�,~Aj��E���XA@�] vRlѩQ���ա�~Y��^��14�x����$T�a�x7Iߪ
i�#�(x�w�h�u��*���Wfw�Nd�0h��*3iG7�m�~�葛i�D�����S��[lN�uM��b�>j����!��P{'aaY'��
�	n�$^с�`<C�#�����d����B���6�A�R�E�Mv�t,��y����t/#X6	��wb暝�8R��5`�ny���C�r��9�-�|�)��Y��<��nos�l����/X{���}�
��08L&�͵v΃��[��9�8Iڮ��9�r^lC�
����*D������^��%�c���P�<���ԫ���-+w�˜��ng���g�'8�EAG��P���!*�7�m�����&а`&K�e��?Q���Ď_�]&" ����&mz�軖���~� RI[tѩo!�w�n��E<�W�V��Y��S'��&���� -��i�ȅyf[X
�O�>�7�nYH�.��jK�=4��	�򒞈O�ԁ�T�:�Nw��A�ɺ@D��r�$t�5��k.z���`H��yD�RP�˻$V�5��v|T�!�J�{Q 87����ծ~67�{g�$��k$�n��5�uk{ѐ��y�d��8�vs��A�r����w����Kh4|�w����%)��MC���:��I<�3�Ԧ��J������gQ��6�Y!/�:���}�,���%�҉�)����������uB��6A%�|���gy`���%�WOy�9v,�6n�}�|~��
wY�D�sh��ut�U���i�Yx^�#�<�S�#�u����ls�0�pA�&�ë�lH��ڵ���jU��c-�K��W��E7����_���t�Sc�(!��z�v^�I�u���]���97>x�U��ϳ�{��x�f��J}i�2����ǢL��(s��n��� 4��h�2�D�E����X^��BE�k�T��W���{���K��W��mc>��g�\C�_�"�@�c�V'�_Q�a��-y��1�\��9֌W��9O�i(��Q�6s҂�#^64����� ����Zu�a���ɣCs�;���γ��@�+$M���t}�5���!~ F �a� �^�ިf2��p���׏��y��@�5��ݨY<bc��)������Sh|�k��\� �->��a�z��0�"������ɽ�#��W�_�	���<p�,��U�z��m���'=W�HI���ATh�U'J4��N(�8C� D��P(���g�L���9	�����T#���R�o6	s�f6�AM&��4��r)!~�3���/�Z�6�a��V~$��Joz�"����s��]tj/��R��{���5�5�|�$�e����Ѫ���*��)�Sj�_N�t�c�ʠn]�G�=F�+1c�2�ZR��$�t'@o|r���qIа]�z�-| ;��E����u�.�bR�$:fq�/�+
|��6�o��j.�"�h�dG���G�U��TɣzF:Y��v�)����5��s�4V��(V�\�,x�^Q���
7r��.�������і�O� c]F��'E)�gV��NH�dYO��7�iriDCH@�'��5������n_�Y�7U])1��}�F:��U���:xyhO���+/��ܥ0�i�^�K�E
ޥ�'��3Z�XY�n�"�NWW	���J����ɱ��\o�yj߾_�D��S<���bw-2���$�T��ڔ�0S��SC�QnSxR��)�[�h]X�U�SD��}��(�G����*b��*�����e�P{����ď�dƬ�c�xS�Rh���x�r'�(#���b�S;�V�\������Q`oN�C�y����.-F��6a _I=z�2�jTHx�QJ�1PCL}�̂��nVB�9��!��D*�R����C$�P��.��G��=(���q`����w�_�����_Eb$?���%�=B�/Ed���D]B���'�n��"�&��L+��5nʏS�F]�T�d����A������H0�&y�=��y�O@���^�,��b2[5���n�>��1�W7Tz ���~�S�:�q��֩�?�G�wp}�/�UQM�	�ԣ�H3�2�l�/�?��2&��g�21���r닖��0�h�#Ŕ�!�F�"���������OU%�"*|Ðd���QRB�5�,!hr@S��,6><[/��kST�3��_>Bx��D����U�]߸I�dٔ�? u_�sj�"e$�҉=l��a�k7��Ǚ�뼫�x����
�� �/���ډ0��3] 5�ɤ���Ƕ�{�k�����nɭ���;�f����'��T�� V^�����tUj{���C������)�>7���cJ�bc�ϲ}E��E���Bڸb`~�S]�� �>;5Kq�/?��9�`z�?�bt����L�K�c�|?t���M�yT]�1W��Hݧ�`}���x��%�kT`����V�5B��t#$Ɔ�� ���|���-�20a��A�2��%�R�{Sf�m���G ׬�JOI�_ϡA���d�+dHS6�O���ɵ�D؀0�u_�߻�o�CD�I���c���
���cb���_s���]�.��Q���������0SL�/�A��3�D���*|�i��AinY~\6=��{�	�+5�I,;v
���X��),q~�9FT�i$9:��A�#*/�<�H��������
��ĎQ� Ä�C�=X�K�A��=�D�T�k�{J��@�S��i���4(�]��<Pt[�d�J�Za��g�C�3,��gs������1�6��G)k���K0V��-�{��&/w
�!���ߊ�����9��8�؊@����d۾��?%BFV��?D�9����S�f,��?���U�^$������՝3�$i~����4��V��
Ľj�'��e���9cv��x`�!��1�:՞~�gK�u#�2%�ga�7�^���5v���=��/I؜�@zv����\ �X�tN�іY����{���f�2
D�){�
m�!ߑ�cǠe7��;�[Qyc:N�ǐ߶;;�����_��A����ÑMS�������,��Niq��L^T�C��"��K@I���Rp����E@��QV� �@�c�������I��
�^q��4��I~�r;-��qK\������D|�I�O=8Y��Ԅ�8����
*hPy�����#�����E��%��}�l��<{�5���
x1�p���E��Fe3�K�6���v wM���J4�8�y	bPب��3��!�ʹPØ�"��g��X��rg���duO�a��l�0ǌ|r��@�7g��-��'�n��|_��~t�ɸ#��xRӀ���5;����Dnem���4ڹ�8��) ^8[y�p�&R0b�ֳ�D�2�``�pZ޷��U�6>i�� �G�.=��t�8� g�v����gH��
����Ю>�Y)�
*��U��H�]�������R$v��or E��D$;����e���f[�:��8����h�ѫ�݉j�zF��L����Z�s�����?�5�"�j��3�kB�
M}�;�5T�&��.DD"�#c$/�1J6�;r�����%�뤰��n���&o��m��~�i�x���R��SY�k&�
�,}�<�]����s��N�`ޖ��#+�� ���1e!� ;g�@��8XXt�7A���w�"OB�����~<{7���[�6���S|+�ۢnf�Q��Iap���Y��?X�RǕ������xm;%ڜ`���X$P�*�ah_������E�z��ÊK����Ir���3�'�h�M!w~k�;pK&=��)l���E~X�t�������Plx�����i���4v~m�wc=����_����S-��qW=rv���2�UE�-z��H�������2����O`�� �o���̹�בo�3�~�����a8�;�3�շ#G��?�gߔM���6���tvҜE &��l��'gE7Wz�MŌ��u�/��v���"�'�^�830�-�$�c��D�����.��O�����tE�^��&+k�}-�3��W�y�l݁*�(���玈Z���vJ�����i�`�(`�ݢDO�ψۛ�!��y��=K����$Td"Kk� ���\��^����J�"�S�=�_?^��M���?�ZF;�����)G���ܭt]���r�ӡu�f��Yf�F��,��%���-�NN���y���ϔ?�E~����~�e>#�e������0&�e�>6\�ZCe��X�,���_@\E�3���e��;5W�)���a���&	1�t���u�$��zW�׹f��䷊�p|pmm?��N��˟ƻo�:�-������i<��՛����m�+~�g��Vv�r- U��z��{�.V.�HU��X5b��ñ�'���4�<ǃ�W��+��V=���[`L
������+F�[�V��n�����I$Hq(�3@@B�:I���%+]�g4�
+-�g��;�}�ʟ�!}w�<��҄_��g�5�m*��9PP� Ol���e�*h�/���~ߍ�A|�]�������2�v�,��ڄ^Z@����1ٕ]��['�\�P?5��-ɩVm,�C}��~�}dq;Pj.ݖ����,J���l��,��!����������0�`66W]I-�.�R��[,�
�9@��١��`�����&��&ڔ���G��f��?�셠ADA�t�f���[,�obۉPܯ�S��zj�5��Y�[�ɸ�,Y��䟯x�%3LEn!��j�PfU�ĨK��\�V̠�3:�	���*�9O�{�{���:���*��M$ﯣ%��_z
Ȗ"�����K�غ
�)3�J��[����7��S\%��ͷ�W� ��3ޘ�Ї��i�H�fԚ� g�ǒt�&O��Ы
VZ4��b���lp�$�X@�E�fU�C�Zk�F��_�*�8�R���6�O�g,wq,�z��VPk�	v�0�ײTV�z�{7��!�`���l�3�*ų҉:5�rlEʊU�-5)���P���J�����ƴ��f]�������2��J��^
H9��>����_%^|X�b�u���iK	.�QWÏ���ѥ��#��`����V=l��t�������Aob�f�ׯc̉��Ӟ���������Y�m"z�!|ڸe} �g�#�g��ՋL�5=�g&ΣP5�GWf���nx��:��_^��3�#`?N�=0��@�ϲ���R�16v�ױ�Z�c�N�?se#����j�&��d9a���E=��.��
qV;�L�+K�N<�6�W�:����������Q�wG{�$�I�jp�-�:ρ���(�|��:Ҏj�W�=���ۜU��6&�pr3%�*(B��n6�Wu1/�&|�&��F�]k+Z��.�n�����=aR��ի���)$���h�[Ҫ��#�6��E�ISQ���b|���8��hOU�T�R<��dh�l�f픾�nZ4��0�����P۱��&k�kP��$���`�(�+c�t�Xf�l�UH�DGuJ�@�'���R�S�S�y�@��`*�6����p��^����)�H�	�d'5��{�f����h?!B\Xm���.����׾+��Xm�7-�$�eA>�/9���U��|�VrCU�����aoq��y�ÅF���{Q3]+�:�L���E^���0�~=o܂̈"f&�>k��,��+�T<�h֬T8#d�ʦ�c���c���_��%���AE_��s]cg��3h�.�yK� zeߤ0�3��kJ7DN��/>�عޝ2�<���Q���.
��^������pS�/s�҂zp�^�<��B�l��ʠX͚4!es�� 馿]e���I��e���1��_��rވ�Jӟ��^"<�����C1�]�N�:?��)g>���T��x����tf���?M�R����}ܶ*{ƺ�b���:Ƿ ��?���e�kf�/�C�|�iA쩞�:ʲ(�@MMn�cP+�,ָ��t^~t��oE�T�lÞA�^�ະ�=��X�47*>�2����ԅ����V���%���FO�&#��ٶoΌ�d���nGI�7ڋ�	�Q���2U%0��7)Л��@D�)�{�!;�}ւx���]6�:���W4�QRG$�!H����� %`��o0@爼��eXG:Dsׄ�:��7O@�zT�B
K7>H�5��U"��L{��^Gd� �/�{c�^G�[�'�Ǳ	.Ѐ)�)O�v�uI��Iq>xT�$�U�+�Q�/��N����y��F��.?�-=��~A�2�Lc�CGg��]�NPn��7��K�<�=/�Y�����Z����5��jnր1fyR	�`�g_Կ����;���k��D�ȖsEk�HXL)�Q
nF��{Df鞌	����@8�P�S�D�c�N��T8�p�$q�Q4��ۆjJ����b7��CG�]0��]��w� �n�R~���3�@����뛔����T�"���o����͇k�s��<L���4��zQ��>3�@��,`'^�,�|�!�MX"���ʫH���D�������3G�݃�r�lU�����Ь��V[@�.�_6�0
m�5�����-g��7��w&\�E�hMw�i���/�_u�+�z�i�v���m#k=8~���a�
�,�3��7�Q�Ȍ�������)�!���:�ۚ.��?C�z���	�?LA~xG|*��+��9!��vX����lp�-�_1�@*�^9l�t�12G���E�/�(�^ީX���߀�rly,٢�	��9ʨ���׳l�����k��k�3nd"�̙�֊߇�^�ѫ�I���#2�����s L�(_��[,��[82�Q,��g�}���k*v���f�Q෤z�&��;�W��4AH��#�/M{k�g�E��ui�&gȘ�w	�4�^zPI/a��e2�j��t��Ecif)�$c�{���m-�a�Ȫ���$���xRhY[5�a��$��d>G��E�$�c�y�ko3�j�e:�	����{�e\m��	3���M�P�^���W&FS� �ь$g3\�����#� ]d���Y�FS��0/�xL%��>ؒ��K�+���1>�)��P`K��T|}�emU��w3�ЂbC	�{���/Ќryu�٦�px=+�e���[׍��GlwZ8����o�n�D$����-z��(�r`��J�|4�uZZg�3Q�ۡk4�ڔy�T ��@2�gU�[9R�У
�����bf��V$���@@�s��5�Y4�����$�&�gDf�3Ƣ�2����o�ڼ�������)���D�����P�4m��}6�>i1�5s�Z���r����jS9��2F�����t��o��e��(À�YS���9����s������L7�B<��`p�=�&/I��Vg�W�������,����ű	�8_��r�)43gٕ��+�#�u,_~��t�`/7���E���9�߻���e���<�ŷ��!�q�y�4�2/^t�ň�.�t(%.�vs�N�����n��OL�Q0��-���U#������^��%ͩ�E�!ZY*�C�G�n,��	z�J�)�H�i�9���m�S:�b�2=P�:.�����,rը��DRnba�U��A�H��s"s�A��[W��.���+���S�#j�b�R�w��L���}�cyw�l�OD���#z/�b=i:دvr��XɎx@���r������uh�<
6q9s\a�ڒwzWV��9Q���V���@f�V��.�Rj���䷧�'�w��;F�~UK�2K�T��r��xw��Ib}��l�mQ�K����,�O-��6��S$����1cX�0�i|���6��|���I�t��U�]?��漡DX_b�O�F��q����K���>~؃ E1�����.��d�^b��`�5Cd~�j�)C`�@�/��7$?)�mɲ�%
N�U�$ko�ld�����Pd�c!�6�@�4�N��=�΢�/��xؗ����.Wh�%l���ѻ	=K'�����:�P�'4�l�KB+���؜��5x�����-_e�S����9��>�"p'^=��k�/�<�n��a����?�2�+~3m��B^�"1U�58��7���C�H���j�h5���?�^r�I�.�Cn}�]/��.��R�8���E�V�5ht�!�O��x���E��^��:ޒ���1;$3��4,���X�h�t�\���[~�&�Gi�V�/9��@�k=�9J3PqH�ӆ�����Y��6���T�t����7���Sk/M��dD �3�X��/�J��+)�2#�� $��b���ȡ�V A^Q|�m��h95 �&47%�<����mcG&�|Z�+���K��/� g�9�-�Np	@�dL)�9����KO�3t�jn2��(m��3q���4�{��}QfHL �N Im�y��P�)\�]��KB�`�Sa�S.}ò�#���H]��g���܆�H~<ϼ}ՊK�	�n�e�́ʭUP��?.>M�5�D�������u'_Y^S��"�x� �k]p����eC��j�"��w�ɢ�#�pZ)�sEq3o������Y�kt��W�W?bI> ����bhN��^�nF��<���;Z��i����A��~�KBއA`�X<p
�!�K���;^��hN5��9m�&h�<o�bӅ��P�B�Z��� ��6i��dF��3����ǖu�G�|�f4~Y��d�q?F���1;���ݚ�������q���Va���ܘ#?�kGo�F�w���;��/�=@����AJ�^�v?�c-�`z�t�tH~M��o����
��,�m�m�6 �"�z'�,� ��\��@��q��'(C�}�*ck�)�e���ڮ�Iܓ4�z}�DZ0;K=J�"��lS��lwj����PO�GB��4|�~�D]7��{3Y��}t����Vk���@��p�`�+X��#4�6�D�������3��{N�*B-U5���{*���8���6��b�U=�s&����~WdX���3�\�)7�w����:^�.<�=[<���]|����%I�嫏s�{i���0N9	�֎�%�y0 �7���mX<����;��N:��I@�e�x�~��BF�&�����V�ޚs�t��Mα�B�腦w'����ԑ�q�5�E<|�U [��A��آ,�ȹ�Ao���Ci!���B��X�'럿�eG���ry��#8��x�F��[�
ܰ����Գ���^ ����_��ɧ���2 ���qNX�p}�E��H��O�t��740`���q{t��A��LX���ɂ�ԏz�OpoL�3d�Qa���fo��j� N����,�GQd�F����8ǭ�Pý'C�ܥ���r�����l2�]�����O�c.cy���aU��ػ�F�ʱ���,~v�k��^��j����u�d)
d4ف�Q!o8�R��O�/��h��-~'L��:N7*��ۀ4c����_IPӳh���1��q�
<�ɦGU���)|�&��D-,�����9���]�|.�3�+�=��[����(�cë_���+&�t�qL����g�3NZ��Q_)Q�Fz$.�'x=%�c���w~�p��1*s�)�h��y,�p��v#`��i�ռ���n���z�N��6he�i����^[z癿����B�E�M��z1
m����qfｼ�,�m��ñ�����;�"4�/�X�Ə�Hb|�
=�O��X�L�0d�?)C������v��@6>��|>�Fɖ��7��I	�}��[�^�(X��{J�k>��֯	UM�2�l�m��uS��&OȥWٌhCZ }d�z�ai�(�6�����(>���l�8\���.m�A2������(��b�V��}c�<�^��~Fu����9��e�F��Q>ʲ]���h�������� r���;�N%�woK�4X��.ф+")T���l�����/��4}�f�.b�ɸC�=7���.BDq�:W�̩$s��I	`E�m��-��}���"(x}�X��E�ߵNZ����h.<N��?C�>�c�-���eV��(�VrE��J\NvH�N�r`xj�.p�Q�g�h�]�.���UQ��u��xp��M2m�r0�Z�n���������PW�����!a��`ī�H�4�S�=�L�u�9D��t�Jf����ԙ2HAD����D��#64�[��1��Hs�s)�|WCRZS����~�N�U�ΒAj*rZ\��&�y�� 3X���nIӟ
d	�Y�� 1���#%���<yf
؁�%�p���/�=�
�[�����=�2����e%Z�G�����Ӏu�L�x���*>�������_j�x��8�/�I�j�u��!^��:���l�/�-EM��v�=A��]���X��i��*~���y�ۧ?\�5�(���l�Αy��8�n�������=�a��۝!���/́�}>_r�oV����F?�R^[�b$ʩ|]�J���Ft\�;&Hj��UǅJN^��(�.�7�G�l��S�},"�nM	w;�O>8�#wD.L���7Α{�5�ל��+�G�����L� �f\��U9	ԏA�n2�T��)��.|����0%���e�ץ��}-��L7cCG[�,Lf�z��zCڅTy��7��q�fD��(Y��zέ�La�u���d�L���r�%���y4���Z?X�RA~}�K��
Ƌ�u_�k��?���C�"X��n��Y�T~Nv�-CM�/�jt��d�����Pv�Y�.��X�M�}��/��b�EJ�b�Y8n�v�?�=j��oS�C��}�
"~w��� �Iq�·���q��;�a���q��墻�|y´��:�.S�oUᄯ89Lڼ	���E��P��AE0%�p!��n�{}#g�)nң`O׷
8)�cE��� =�^2�4�%��k���o�Q
Nu?&� D�fvë��,�F��Ї�H): 1\VK4�ޜ�Ie�'�k��k�i�9����]��JA���Z+dq�s�o���7�Zun͍yK2�����K������DzϘ#��</��rOe�k��b$5B��.,x]�<�R<�����{�L��Х�������}�D��C�2��7ʾ[bT�cH_S��y�ekI1�)�Mp481��&F �ƥ<Q�=�
�z������{i�e�c>s�#6�\̺��4q��Nƶ�kE��c�%l���j�~�k'��K�.d�p�2��	���P���
\9S����<�d�\��m�G>����Qg�ܶ=�O�	2�S��de�%C��z(�L��������a���w��U��5�\�	��p��[���,y)�^���.��B��˙m\{H��%`�.�t�
����K`[��*Y�8|�D�6,JZ�Jo�����j|}��j��`.���X.,;3ɬ��M����6N�?5�s��y���I�"b,�R��Ǜn�Q�Y��/�q�<���h�̳�<h�E�Y'�ql���P_�0۱�iuL���k+gC^9e��kt|~�6���@n���K����f�C�F<��LG���H?�����b�wF�
��s�Ƥ���<1���?������˭^)^	K�RGZzrk��J�j�����������R��z�[�埜�>�E�Os.�w�W�լ�e6K3O���I�Ih6D��]JEa.&�Ԝ����i����F��p֍�1B���_������!sf�,Aܰ�,�ŹW����(��f��k0�.�!�VOP9���ݼS1`q�|]�8E]��*�X�UU��M�  �t�{���$? kq���\�`�uq�}S@ŭLv&(qș�"���隃K���Ϊ��B��p1���eқ��EjH�U'�Pc%����~8^�s9��<����x�'�׼$4�JXD�T/![R��.V��m�?�E-�\Hn|J�c=j�l�K��F~R�_��aS��	�G��Om���[��'��)�����}� �X�"�P�	+�6��`+@@U0���{�rtʚn39��O�{w���Q�l�FZq,omb�|�t�@x^����KK��8����q�W����]� T�ZO��> i�|���}BWkj8b�sC��G�R�QZ3J�i+j^�|�3op��/�Q�'�̖C����S�%[��:�oF#D�KD����W%K<�wޞO���㹼��߾zF(٤ʳA���?�7U������a��
��O��y�k��*�����Y����\��j&��[�u�	=t����/Uʯ�� ��C��@$�����`��Hx�� ��&�6�/=�_Mr�+b�w( ��d�D5"5�t%��zߗ�$�m�2KO���@�8>\�R�{z�8���͏���z��ɟ
hKr~ES%�3����n;ՆB1���\�[� �mn��8���ڡp#�vZ������G�w? �$��4׌l��@t<�̝�p΍��VM���#Wl���L������ʸK|oz�
tp~���U5��g�4� �Z�F8�J���=����~[B(����d����Ϟ��N}�/��[jx��^������K_���lb���'�Ic�Jx�*�zZ�ϻr�������Ȓ<��5J�϶QO���:���>�%D.G��@6���Om�m�:g��bC{&�q�W�p��U/WV4�|=�ͳ랢P�n��'x.��rJ��+���o�'6:����|I�,�:�������2	�(-�l�SsK�
��Q�>��v*�W�)\�{X��h|�����,�J\�Ҫ(ܜ�x���� ����W_X�	���;����*��N������|�U�������0�v������w�u�|	����->eu�yɱw��}юJV3����DX�-I98@{+�����My/G����gju��ߋ<������-<p�fw�z$���s��B�'2Hz�[#��W?S�����!X�Ӹ��0���B|��&�A���=_g��N���Id��G�6OW�X�Z:�+P�R3-]����q�=GZ��o�yA	cnv���x�o�y�N�g�$M�^�����z�*=��ja�.!���?�+{[�E4��Z�Utb|n��ԼOd�jגT(��*[Ol����|���ek��#mi8b2�����U��V��KM$���
���7�{]���bt�c�T^�Q6�>�oV�I(���g@�<�
�b?���+ ��.�yzӊAF�8���� *�t�w;�^*�hw����q�o�
C�^v�D.r�}Zd0`��ƽ�b��l�}>��{G���>�TH�Xa����wn�oWa�q�;,PM ;_8�+!/���ޯ��+n�{�ΒH]�cs�x&}��� m�HuX�	��1˨QEs7̖N���Y�!��ۓ�.�!L���k�R��_;����� ���Pi#V�\��Cnds!��q�S���0��2QU�BцL���
��[E�B��n�E��)����/ǤR	T�	l�PL��F���/� JxLY�5.5���|C�U��RlwR3�A��7F�7ے�����L���Ԧ��F����[�3A���P��Qڶ#��BNZI��2>�Ѣ�d�5�w��
��_��8�R>.��ᖂ}��U�R�˔�D�u_�Ä�l��u2~>������k�wkS�V�.��L�S��/�lq�{3�&��5"qR�cQtުCMFRǉyN�bS����8�<��*���h?m�'���R�ȳ굉ZZ��&��È�%/�$����F_�#�sc$vΗ(�S�t��-�^;C��B?�����LMnr��D�Pz#��*.fJNT�:e�i9��/�K:�6c .zؚ�}é%x�)�Հ����s����@J�gCOH���o6��}���oC�A��sZ�v�Ff��(��O��^�Q�����Ϛe�/����3:^ti��]�,#C���T�($AS��Vw���|�j���1+��yt����fa�o��/�F&�7D����C�vX�!T�&]������D��B�������|x���-#39=�/���N��n�pܝ#��4����ev�|�R)J��b��Kh��LXcN&�:lz�w��db��L�p�[�3Q���	���Z�ڒ�qs�ruR�*�������rQ�=��!�����E�j������0�|F������z@S,rr�������Ia+��s�/uQRC[��;�t}
�Y��b;��:ǃeA��>��}F2p@�uJ<�t��`�b�ڌe����F~)m����sH��[�p)�9���M�ؾ���ۚ�ͅ�g���$�s��s.�eO���M��6N�L�5j��أ���������k;2�N*Ok�m����O�>3�م���6�
��f(�i�@(O>~��#��%�2!u樤ht�wX��[�
��[	G ��j'wB{_T	ܐ����j��R��e趼�w���M����b�9�xM\��`R1 lt�[� ��[�%���Q9��"$���t9���M�zIF��c����'������I�T�-�EenCB�6�g�+��R>
��Ѳo:�P�;�GMvʤ5��!��#�9i2�TKL�rR�������z��A�
��b�F��{�W�Z��>M��Eh4ǯ�:N�Tp�k�)��v��x���s@��B��5~�0w|��N&#X�,��*Z���Þ'���OJ7]��)n��^�4�dᐞJucT��?"S���$&�@��o�I��D�)w�d���W�9@�g�Dl>�3ß��e�zFi�{ z<��T��Qx�s�E�F�
�nt��Wm����
69����(��=U�����ɣfA9� �����H�7q��P�qy� ]��2�����`�C3ol�C0���Wm�c[�N_ gU�	�}ݕR��~�،�������*!+s,؉|�P�<��{'n��:��f/Z�gu9����(b��j�I��Z�J��D_�*m�������7��+e-���^�ŵ$�=�d��`oQ��P�>7�?��Q���6޲���fhPf�f_v��s'T��T��G�a������k��(����s1o�j�FI��PMfb�	*��r��F�"C��>>R9�\�V��������=R��(M{�X��\`;��/�Ŕ�
.!Gy����Ph II+���2��#UU�d�^.펚.�s�mr�D�S�o�-���i�w�N�EXq�m��q�0K;י�\�5������/_�z�-#�X�_c`W�¡�-��O`��r_�h
��6]�
0�o�٥�Tյ4tkӁ��y�n�(��%+,^�[�|-�}P7R��2����Q�d*��tyt�z2y�޺L�2�*�0�ǵ� [Y�Fs���_;Q��ꪚG���\����,A1���n���@8֢U̍H׎�Ø�e�MG;��6�=$�;H��Sl;��B��8�S��My�g��*lH���\*�q����������3�k7svT��x�;n$]�RF3��s<�ew���b��V%�s���� 'F��K&�!��gа��@g�O��l�u���a
��ԇL��S<�͐^*v�a�f�<}+W���ʜi��b�x:V���_��0��;z޿�	s�>4?p�S��S�l�;�5Rvx�3%ǽ�HZNΕp@L����	 |��l��Duz�%wg/�����p���K�u����FME.���Om�x�Cz׵����y4x�y����h��,��{Mȓ+Q͖�j���ɍR�^�V��-5D��pÉ�8��s��o:�W]Z+��P��ƭ;�(�2q �Wny�@^�%��Q���M����J�� �;r�׵RXR��>v�ۅIK��^�;�k�����Y�ȣ�����J������zǌ��ސ�){�9��*X�7�UC|��xﾧ�g<�/���]Ჺ&�����f\��\��#
��p����{�h7&���Ի 5Z��@[�ja�HQ�'��D.�!�Ty�ds��W1ـ c@RƘ��?h���#H=��$�st�Z��� �֥�0�Ъr�S ���=��g�̜�e�"������H�w���$@��;
�E�<�S�$]g��t)7J3�и�n*�	yE����aZ7�S�n%�4��_䃻	a���ߋ�� �˵U��"��7�S�ЛD䰇���ٮ��9w����J�c9Z~�7[��F�$�o�~������IC�>�<�����Q�P��Nj��0!E,0UNpF"B��`�8���j�|�͢cܚ��y�Y�[l"��t?���O⚴n����&������P�  �g`��
+=G��=Ӟ/M��ʕ���1�Kʚ����2���55\���xC��pmaoA3�{4�VG�:��\J�K?e0:��ˁ�S��7��ۻ�t	�\R���)��6H�a��#�Ea@��c�'�p/2f��:Nl���YW�*3�Z�O��ffR ��hqw�����0Z��j��Z_d��q���c,ƈ��G��x<Ӎ�a��5�9.���>n�&�u?��jh�<�hJ��`�0HA�"}�#@j�Dq{�ef��l\Q����W](d�?��$�\�Qd�W`�eο��6-\DH��Y�i� `tSg�J>3?�)�i��� %z�P�hK*n�"�U1��y,KD�q�5@;,f!&�ZX�)�P�r��Hs�47���q���:�(�e�~8 Ϙ�5��W�M�g�!�Y��X~ٽv������/�SX倲k��Z�8V�a�MKEf�_�QO1LɎ����zV��eCT�H0E6����#?�lH���\�0�7=.K�W�P�����#� Q���ew�R���	�Ij�y��O=�.9��m��Ԯ�A���d1��T����ڡy�f���%���{P���S{b�=h?�y�x���Y"����?#7I%��MJj����U��#?����6�Fcϋ/+I��+��@���|��e�d�Sxs��G(:TprG]�9������V����U o��#�	)S_��HK5�J�A�6�$,v�����9�<=�N�I�i�W3f�%�p�0��;���<O��_����ҴVPK{R�Q��Ā Y��)��b �!'���d��h΍�ƑR��Ɓ�16w�-<��m�����4�沸���j�CZ��i�R+��Y^ܠqG�36�uܷ��	�|�jk0��Gv,v��pj��	+E�[&���*�4M�/;��_���&OMi1��qUT��ƨ���ͱ�QP��e�c��{��f�H���ao���wq��*�����>��6>�9��nw��C�+v~����D��}���hG��r0���=6Oq�meԸ$t0.����ˡ�FtZpM�8dK�I���-F�9=x1 z��P��%�g`)H��X��UD�?�㌰��9!�'$��T�;˶�~��PЉ���x9����)�b:�4���L��y�Li1�Uk�$D�3�r0�%=:���W5�h]Ԝs�7��wu���o�mt�mZ?��N��m��ĥTA�2�z���r�����{zZ�|e�Ȱ�!������Z�~f����]_3��\�V$�	h�A!*���Z�p�UR�I��؆��gGi��ηW8_-��M��Ž��w�%2��A������Pr��L�T��x��hŌ[S^�:����fp�����i���^�|t�~
��و�ǚO�D�Tx�AZ_A˸�~���@n����C����Y�"B�5 ]�gNx��G8G$U�V0����ܢl��ì��K�=G��>e��M�^��̤�ܴ��s����7���,���o.>����t4�����n�(��=K�P�cy�������fT���`����2)86<�4����]W�e�
��k��{��g	E��D,O>p� �9Z�-T�
�s`c��zX����h�i�6� X8�
�lmլ��zDjš��ף� ��T�=�|�# �{�-��k"�!�x1��ݞR�sq��h-�X����nk��Ք�.��ɫ�TBAM+���z·���x\Q��Ӳ�:zq�0�����\�؃�ZsHjJ,0�ŋs����!�On�O^��G��H�p)qڌR � ��? ���G��2��HP��wsV��Ǧ}	+������!�t�\�>V����k9�d�ҙ54�Gm1؂NI*����m� �L����0�i��4�4Θ�a� 7�ǈ0ŧ0��)5������p�bޘ�W+=�����\����t�B�pk��K����JBt���N�j#Q�r����J!�?����))y�Z%����4���N��d���cuj�*Hv-Wl������L�r���fԌV�o�c�˽�ClT��$�dY^xNnejb�re0en�u�6�X�7/5�Ͷ�eĐS�5A�NTCA�o�bI�bi>$U��!V���MUG��d8߅U�	���3��[�s�yn����dUOk������� �w���4'���A��b橓7���{���*ώB`����4l����A?^�t�QX����,��v�a,
{�<Ζ�%�5гE\"e��?�0켽i������|�d�w�_&�`�`b����;M4%���	��kA��=�����q����-�?2������Y&��Q�������6����ވ@�?��l��R9L��Jacj��_q�6�:���M��q-�(m��g�}n4k�H,i6�ߙ����R��'����|�⑆���tj�]��w���Z����?����G{#����5��EY๪�����H�y��ф�3��I#w��_;�O�>b?����U}g\��68��[Ç4���ܶ�ڹ'�.�C���c\V��<|4D:SO��{$��k��!D׉�[�xo&�4ot5���Y���.��5�i,�5��/W��$)\Ls��b�/�!�"�����oeQ���|C�L���c���o�O����^�7\��b�z��o�:�3�Kj���懠)���+�5`�N�FT��0U\VB��$y�MD���n�&��c�������ա1'7i5	�h�(��$�c�5g!�A�u��0?�fx�ެ��vƄ���VxUS�bu���z�#oЏy����n$���e�-fI%��)(p���_��{� ���z�8d:�Z�~�L��/^��?��mo���#Y�/�ѳ�����F>�s��[�!3(��ĳࠍR/[�T�}�@���0�Fy��m�+��Hl>�
�$�d9����*��( ���<s�E@.��]ΈH_"��g]�[�m�az�D�3r�>~�$�>����CJ��ew�m�V|���� �顭N�ԋ����u�>��/�P�`�='@hqVa+/:9ǳ�$^�p\d����3�cjzٟ��^�Å%�pXH�u�q����&��]���#6�`4n�qs�C���S���r�=��Ƥ���w���ʦw��dD��?�=�G�^Ii!%gckX�(W!��ˎ-��ԬHq�CTv\d[���7B��C��5�)cO)*�_��x{���i�����(�~� ����iٵ,�lyn2u-F-�r5������M�"�g�(h�Ԥ�8�v�6;s���}�o��w"8^o�����y#'�?�8�Z��E��u^�uT�O;�
�F'^2P�Ab.9��AE�iw1���C;F�b32�긐]|"����NEs��8��/��pU�ͥ�K:�!3��T�Z�You�0�	$p-#�țV�o9<�Cb�LM�sӼ��TH��
��<���h����;��K�dQ(O���%0sf Y�	3���+�\�v�g���/%[c��h���B��/{I/��E(ش3*�q%���M�35��X�
ߣ^O_�~��/(4m�0��dr3����yɔ�gB5u�A��@EYd���`=���G�·+�Рj�N4�}��2wudn��R��Mk>�����a~��y;^�lR�t}8��p MXwܸ��	�}I������j�k�bb,��o�Ic��6��t�Pñ�JuT���aV��m��J���a*K��_�M�l�4�)ycq�T�$3��$�+�-��ӿL�Wƥg�~/��K1))�)t�S�+k�X*�³U�Wb4E�
�5�%��/Y��TA>�̀Ir(.�bO~��PSp�'�d�o�g�H'ݳ���HJ�?�Peߡ�̟�K>mhV[ZJ���36�%8\"��S_s��f(��d��'��^���������˽���<��|$�9�����N������FUP��UB�
�EaB���F6�/B~�n8b]/t0}'@wWb��j��-��Z���[��6��r�n= �5Ǜ�M�  ^��f�-������j��?�F8�L�%ER�ߐ�܇�2#�SY���l�/�cJd��y��x��2n�N�5�HI:*��11=����E"[��	f�n]&E8���_*kamyՂ�>���:�)bW�n��ܴ����V�}�|v�\��ׄ�d�+�V�u[���[�q�2��<�߇��g+��l��9'U���?pr�#�D��:FJa�f�Q<�|L8��g	hp.��۷���y,u�8�K�� mђ����PT�R�4�2e�VI�9p��W� g�@.��xH�"u�&߄�e��?e&3�@�7�:������]����A	c/b�����iO����M/iARg�"ڦr
��ρ:�N�E�9����g!x|Y�����F��=շ��5z��ɽ�՜ר&�jE��qCG˗��F2�oa7�nU�QXUNJt��?�5�����|�5�pL��^;E��mBi/e�0�4�6����X����.͌���-��.�m�c��9�%$��lc��}�{-���d�d���u��=��B��/<zn�N�3�[8����LZ�Cw�Ȱ
�^-���N`�=������E�Is�5���'w7zrD&̒�к�|��Iʫl�.�N�l�9�˯�&G8�Y�Mm��:�W�����I��D3���iG耓�6��)rQ-��Ӡ ��C��<@�[lZ��s[��t,���[�>) (lri�)�V�c�YC��%x�YDZ,��_1���|m��N6���Y+\`O6�v|��!����^��	�_�t�f�,����Rlƶ��s�Wέ;4�u���<N{;2��6-�O������9o|�l	��*0(ַ�|HyB����{I'�e9~@�9YtGdW̗�h.�u��չ1�f묋��̭���t@�H��@?kk�T 	��y?�a��hs�� ��+-�-kH���76�;��]�����
 R�-]�ȧ����,v��&��*V�ӷT�$�΂$wh�ε��3��𾊣O��%u����������c�fd���cC�B�7t�>�@W_���d�[[]�+Gork���}	�&�����	�e${gz�cH��WNmܾ���O��r��2�c$��Z��9���R��=�&�$�.���LW�g��V�K�q7�\3m�`��	�E�"�:�����-Nup�1���_��%��?� ��6�� !�A�h�B\�,5%���9	+�}��{g,�� %|xE�1�2l,JkZ��)�}���}xtwY��qV٧���f�ԁJ�m��\	�F=$���"��BlU���:q

�%�wJ��3"�'f&dIw��;��Kp��8u�4�g4_��Q�����.)�d��QB���������b�~"٤ޫ��O����<��Ú�i�"{�n�f8ܞ�{T�h��;KA�t�3?��5��HA�3J�7�(� Q;����?
<���97W�qf��M�Q��N�i+���/6V������Ď�H����H���tʔ+^�ެ���?�\�0i@��P*/dK�U���'K�N�A��O���7�W�a+Fcu씑q�;��ݸ�XKTFLY�ӫ�Ő8l����=#&fe�0��G��t������{�"`Ə�:� >h�갂b0B�'7���0���Nw�=���?���+��<�A����4�yǙ�v&���(�����?L��Vq�UDJ���A��H3ž�������������TGnc�Ƞ�j~Rm ��� �uu�kE�ѿ�������|0�8LD%�	��:o8����]A)��-d�+Ty��L�ј��.�ƵP�,��;nQ ��H�����:n`܃M>�X��Ը��2�QuI�tl%�PYm��E��T���ő�y��ABo���YE\��.6�"֊�0E��z�_�����o%�8�'=V����%�bߨI@�:���b5�<��(���HF�!���/��[{�:��}l�r��TV/�nV,��ja�EO���V(�;$'h�5���vu�j�"��:cd:��C�]�4�=Y`�Ԓ��pp�ſ��b�c��g�����`浇_E�c/�lɞ�l���~Y���D�,]zx5�^���,����6m�;�5Z���"����[�D�H�,��Q�`��EP%�Ѝ?�p� �VԜ�\�x��<�MY��Xˠ�$�͟ F�����6���m�S0�����O����L4�ˈ�_q.�U7����O�&h!"���v���i#�qT.�:i��'v9k�yrI�yp�h�c�ͨ�`�����6r�f��pm����:����8X�jO���H<EV��Х��S�J��J��~�I�#
���d~02�֐{�zi+�tm�K����n�#�TX�P~6<�}j]m�I}�A��10(�J�R���-㬸����C��]�:(�8� M���v]� m�ߒ�f����R#�i�! �������
&�=��q�^"p��jt�9ψOS"���y��>E�q�ūaea1� %�̠We�Ψ��$���֖���忾J�������@���>Y�v�(��X�I t���*9'T2xE��}`b1s_ڍ!ʬ��l���g����~W��c�H����IPpe�v(+Wc�������Y���&�]��t��<�dz�M=c�n
3���f��J�G�X���G�3κꚟW	`�Ƒ��^�/b4J��g�c/Ȯ#�9K�}CC	]��@ʣfܻ���d�����K�\�9Vj��Fp���c����v�zԛd�D������y���'���%u�V��&�����������OԪOn�.ݼ��x��I;�M3��PD��_�y�W��;|LqG^�W�6Ԃ+[����	Ljk�I]"�1�$N����)�X��=�������H���Z
<�+w�@D�Xk�U�g�L��$�����um��]oYlFc�d�ڨ���_�(<��E��y�r��t���Ň�a�U�p�k.�mW~��H���l��X{%�9;�O[��V�DԜɄ6P{� �>�SPS��h�54<���H��c��XOI���d��maؐ�2R�A�Q��s׃�b��[���H��Q)I����9�pS�M��+����r~mp���@/�)V�fl�Ok���Gֱ)����f��#(9":���E{��Z�
i�uk��L�YD�!.�b��:}�<�>SB
�0&+�[t��Fg7���&O�x�8�V���`�5��Y�:A����oUh�3�v0��<^�a��*PSc�w4��C]�0�gLw��-|�^t0�ק���RG�J�M�� �4��~��Q��4d��L���U��N��,^��Gs�ۿ����x�����"N��_2��rl5���%-������X�c�=�a�);��|E!�z��4���(��ZZ&9�dS{�;���lr�����g�-���܏�R��|��^\y�j�k��[1�G'�{�Pލ���_4T�-��jw͋e�I���,/����2a�"�n:P�$�ߝ�|���D�����O�&wzx�]g�s=�eѳ�%���Om�
9\�)�J4�ި)_TCf�l\ǃ�f�* t j!-
�0qA@�Ƃ����Y�8[�o��#�������Nbؽ��Χ�Yu��������cY
�e7o���:��#Q�j��B�� ,���IA3����.�=F(K����Jx7��e�����(t�2vX*"xF_�r���jj���C"J�^���;A����|2�dQ�������.�x�=���A=��z��}�aRC���5p��ـPsn�>I�I��j��X��*@����@�0G�a0::�v����M��_�Ľ��1��]�d����!��n�7Lb	�Xc8�관���J���&�a�;���`#�gB@��wV���i��-�|���'� 0
��Յ�W�Fȏ��|�"�K)j������µ�7r}L�
鯧�@�B٥-�6�'�e��ͦ>���n�?�zL�7���/��[���v4�3 ���J	j牿�8n��8,lP�c_��p�Y��Wc�1����D�*Nޝ~Zx)-��0;�8?�v�p����.�c�iIh
�? ���$�8?��l  �e�Y�p�`
��c��>�����V��c�~�O���P,5Ic�9�nf�s������.��]Z���hԀ�n5��R��ul�Q5s�E��-q`�޸�^�b%���I�z�8}=��g`�K�����ƚ�z��?nTSO�M*0=���yXƮ�?낤E򀤙���V�7�A�[>�:K�@�=�VG�+��5����}�l䠠�V�v^��.ٱ�XږRD�	�uP�ېS�y�P}3�h4jG� �|�{.!�E�.��_���O����4Kh�>��|6�z=AF���T��`)n���J4GH�[�=]PV��(���-��j�/�Q+��4��{}�>��vr&H�UsÖ<"7�>Gv��k�r�;6��4,8�V���H�t4�)�S�nc_�	�:N�l�	%�d��<���X�L2����+&�zՔ�5QZ�X���ڀP=ǹ\��ЅBeRÍWI�)��|���'��*���pHV�����O^+�*|s"$�w��|����Ќ�����B�J�? ��5����1f��߀:�D�>�OZ�u��qjª��
L�D��Y�⵺��	ba`0�|�����O����iLgx�
1��[��H��ٟv��Zwn5�?�W��7{Wy�-=�&�9�>�o|VH��p2�����	�b>�r�*k�}��ѧ tp���p��Mǘl*��!���NJ��-F �Ty�^�[j�% �#\F?�N<a ��&�d����6�ڣy���J����nn:��6�|zWZ&v�:?�6
�M���܊�Ya��Z����?M��Q��"��U���,�����Z�昝�����Z��d[�R%Ē�X�(G�}ZT�� sL����]c��3| Η�y�yNXL��)��x,>쁬=�q�\��z:se7�ɯX���T0�Ҁ�`�{��ߛ�b�6���Ó�-��o��}�3��ŁlE,J�0��;>�&S�-ΦY�\Ӑ�xC�8b�����(��ryǂ=`�4*���w��5s��p� S��~rh��/by_i�FOC���rm;Hyqw�w`�AZG
�#h�#��ƪ��̅Ν���dԷQ
]���<\�[]��}��b�����3H4�%�F�vc�U3ņ�x�O�Dˡ�lж���Qm�>Tw ����ԣ�qQ�����奃m��}KҘ�a��S���8M�Zw�����n��PsJeٱE+k�}�K������6ҹ��d�ٹ��<����6�E0��T�,=$>�C�K��|�f!�����Vu?�8�v��t&��a�{$�X�L�f]׫��iui����^M�A�(e�=���r��Yz9��\���.q�B`@4iŪ�̬��"L�?���j{�+z0U,i���8���B
�A�������P��.�זE�5�Τ��͡4���К�4-�	r��0��R!��Bn���!BR��>����n�Y�._��+O�1�?x���_�fl��@�+h@��f���fF��^�F·���6�r�qUb��7��@+\���PV��l𲒼�7&q����C��|�J�w ���v���o"R��h�:�JѹI�Z��4��˭�	���)#�r)_ی,��	¯�H���5����%gt�u:dѡ}/S�,�)��]������vK}+�V���st��/�'��h� ��=L�p
g��4�L�uW��㩼�=xCcOkp�7�P?&��(��C)rJ�,t]�2N͌�5������2۞�'��;��_��a�羂P91���װ'�CK���2T�0�2�����pd���g{��"BY��8��J��kMlA=����a�aK�"<4H��uB�`���esN�k����V��aJ(2�$l�E#�V|�[�ޤ[��eb\0M�=pt��`'7T�k�zÑ���v@�;���@z.��/+�>��{�S�u��߁����5�s��^�S;����_�D+V �A/[f�oR.�7@�xʺVǘ�c �u%��O���m�?�fIs2�(}Fj�U�F�>N�`��@	�eyo��*��ɼ��bs�_qtr�[N.��;�'��7�R�ʖ��Zi���i��E��=�-Y{�bʖI ��Ł\F�_aq�y]�c@Q�?�̮A�L�Vc)¹��l|<g7�T�V!�:k���°s/ڢ͌Zy��B4"�;��^׎&�+�O��s8'|�Zr��$��G���(|4D���
�Z��hҎf��m�	k��ȾM�����QR�ﴠG�,�0!E�IqM��+��||ļ3�%�tFY���r�=������J���O��]Ȱ2�!�(�(?�13�����ښ���P��eB���q��'�N��K�t����h�Cgi�3����s:��B�0z�K}�>E����(�L�1��d�@��=z�V�ߵ�Z	�F��5����
��˅O��(����]g����m��lJ|j�%9�8ً�ؤ"����0����,�»m9�M�^�zv&�=,�K�]��W7+Nj{-���ă;C���;'�y�3b�0�ѻ��u��q��X���N���1�G�0Ǿ����/;�R��xܽ]����pG
�o�4���q��\*���� Un���1F�+�Q��H"�:���*���v�D�SsW�#�e0,�.�IzS��-�N��Uӵ�����7]��Ow�dW��ȡڛ���x��2���%KQ(�0&k;�"��b��E��w��P��� y��H�O�U���#�u�mYл�~��6�3���*�M#��!X�Q����`�ȴ�	�M�����x�@R�ߊR~\�e�������˯�G�1�"a٠v�h��7�����8�顝���ljp(q4�� '��Q�E�+j��;�ͺ>g��ǚ�LN*�˼I�i�R�+��!��_o�ɣ6g�cxQ4{p�H�x���M��f!�lt((�ҕ��Y�k�}�F��b���AM��s�({���-�0�w)Ќη�e��ĸ+����ʤ�`{�yI�8����JrH�:��������)�P�\�u	.[��S#��iKk`p���FY�����N�:psh!�}\��L�G;\�F|^��u_+N��5�9nA�w��՛�s����X������5ٯ�OW��d(�C����ð���}�f�Sai�'��"�#7!����F�Z�U��%I|�A���b̡82hƼ��&Z��)�)qx����GD�OG���zӠ#������ɴ&���B�&80��+[��n�G��s���%ײ?4"	2$��
��OE��m~c>bx�ŃD	I���_P.F�'�)Nn�y�B`�Ε��W�|���[\]s�V�4��5�+��� �u�=.��*N��!-Y��砑�x8t���s��<�귿ɘw���8���yX�����wl٢���Vj��d8ў�����h��(�v�>��η�G�ʎ���H,����W��֨{��=�>��d��J�*�
������Â�*F.9@�68���0�B�N,!�*{D�yټ�T=�X{-f����t03~��K��Fr:adl�1�j�4��W�X~����o���U�Z����{��8 �	�ܹ|��&Q�nDU�3���%rg�q$5����/��������G3�/��\���0h(8
�R-_Fh�x���F@U�E\f�)	�K1�$
ub��R]S�?�R6
�2
�� �)�5Sl~�Na�/G.��ئW��TR��Z����lƇ�+�'7�"�Kb�4��Ce5 �cR��Ҭ�p����|��z�lzs�ǽ&cD�L��`��9!H^�����9K��1��ڬ.L!�]	��kqI[��>-Ƚ{FS�R�IU1-_�N�"xr�ui�w����^DvTʯ�����9Hz��r��S�d���k�S?�֋�7<d�؝��z�CQ��7�W���$0�����}H����̔�ݑ>�2�4K����/c�:���>N1��N��I��)�77��MCM1��j���q���m��XKo57d|�r�t͎OKִ�9�
ւtO��.?͢�TfL�t+��{���������K>)1*����V
J��J���H� g���&H��.k�͙#��x(�H��E�,8�èd�^M���ܐ��������!4�M��6��ý=������7�c���ǆ8��ؙY��#���sw���55ق��5���_�'z������>rBX��[��(��Ӆ+�G�?O�W�
�Ir���8S�&�Cx�.�g������S����-@�ʩ�{������n�A��:�BZ�N`|Hh�(r�\ˊ9��&a%/?�t�ĝR�j���Ǯ��ȳ�ɀġ/|�M� �Rwf�yƧ\���+O'���h��q��8D�	+�4�Z�<�1�*��l(��Len����i�w�v=���a^c?��ࠒ�"���`��I'�y�QI�����3�0�b��7�ν0> �Ur��*5��(:->EhE�^�<��KC����`p�,[�,�pD�$�����1o͍��=vr-�A�{A,��z��f�)���%�|S�[-}���rF��3�L���|�4��������=�N����f���-��d�
��؍!�j�I����Z� ^r���^�!x�O��z�����zɏiݙk��R����7Ѡ��E����e�� ���?=t���������"�$H��ej����sd��S)�^��:tާ� >Pǻ�}.��Ga���#�������t
�m��N��6�w����la�p�$K�Lj�_�a"�WHC�a����������a���T��-�̍���R�?͖kB��9����D)O�e(f!`Sgu������HNB>�CY`0���#T�FYܛ�
�,��6�͔i�!��:�2�����N_���1����)ö:�#IQ�3�ݿ&���`��)I�5;E��X9mu��-���O�d�J�j!�� #6�p�3���ޤȳ�	q����g���4?���
�3\ŵC����������\'H7�){15��!������ꂆYq��/��5�-�;��7��� ���%oϷ<��p$x�1�$\E~c����a�;VZr"�cm�r��������l�t9�eX�W,��I��`{�N����l��)=ѵ�1cD?6~U!;_>F~3P���1$�Nb���ot��}{!�;8�I*L��3�rTK��\"�:M"�x$"����ݚ͉�mbj�j.��YK�PXUp �@���{g�R���s���c��vU	��[�H��A�i����<�Dt߫���D����_�"�鉻(L��"@�s�sʢ����/� ��\�}�R�F��+ͽ
ъ�6�i�S��U})���>B�C{�p��}YZz���[w.[PVTd��ܤ�;�ڳ4E'o��UN
)��<h�&�v�V
����-VM��M�=�/e['���s�LG'���S�֐I��yY��mG���u:*������>�'����
b ��XK�'�u���2�Pǰ�����h��`�VBŤ��i�G��h�`�fm�9��#r|�?=���� ������s�Հe�r\��2��μo����GVE���P�\�r����UW��/sM���KL4��YP{�+}e���s��1w)�D�^._�t\����Q�Q�Y6GU���e3����>���+I*>�p��X�Յf㠳�Y	�n��՜�v����շ�ݷX0�]�q]��ʰ&�B��	z=+�~t����޴CB��s������R	X�W�"/>�J�����4IT�vOǑ��q�B��:�Tњp��m|w��s���V&��	�-��XZ}�v޷��B��:0��/�px,�>�ሶ�;V�IW\)�q.cwǥ���!��AA��"}5'��R�Ճ�ju �?
�Λx6�a�Ug&ڟ��V�����v�3§��gTN�F7Jl��F�y����4^��'�|���R(��.ѻ�֘��=���\��kۜ7��۴zɒ�*dY��A��e��3�j����B�.	O&]��p�2�J��K+'�=;���:�{.�'C�!.1�rZc\;S9�{}u��j�EY�m�*�Z�
8�{��ŁZ|/�(|	��ǜ��vCL���=�H"��q�6'��
�x��q�K��xay�KG_�bM����I�]1��	Or��B�L���u�xb{m��j��Ϧaf�+N��\���TVB��������u 1�_�g<%�ϱ���;����T>&�CO����P��r�*��L7MN��>a�$
z�f�E&�e>N�}�сmG��T�Tl[��տ�x�KB�=�^TR�x=�9�2�톇��"a��#�����e��P��-ZF���Lx@���Zb0X����#X�CU5g"�P��1��q�|�bG����e��Tg:��o��-N/�a'����u�|d����ۚ���. ��HQ��=��ˁ�z��c~@�}9s����x�-����x'����y��y)�;�;,���䯺gj #��j5��
��6�w)}([�4�9�nX��>�(��h~Ԝ t�O�b�0��6Ɩ����;�����d�^Ⱦ���ն3�5��]�5�NCOu�'�Ni�
�`L�]k��g��%|0A:Mu))�����7���&XK%?f��5s����� !�6=j8�d�-E�k⻟p��tX��V�9�(Y:���Q��@O�ڊe���8�U߈8DF�t�_s^�{8M*fce�P��D�d��ɢ��F!�C9n�XH�#�����3N��i��3�9��������.�ed�!�j��������J�~EƓ6M��+��ݰ���C�zS�u;*pL��gL�E�<�\*�@��x<��#x�8(w{')��8�=�����|:�4V���#�n`�D��1�ŬA5��2oy�����R���ԝ��?��WE6����� ��BcQI���K�� G
����xd�-��M�߾��TA�$7i�*����)&-�^����P�R �O�pa�:�]����BNE�9�.�Q�u�;vŹ�����0��Q[;�dT��X0ntd��1��Pm�ɉ<��Ȥ����H$�|6�gb?�¢(J��v�����0��:Yj5=7bfgs,�*z�J��g�	��#�ha�#�Ⴑ9�E*k��hR�	JRԲpOuܥ[�L}���J�C ���x=POvӋ�ٴ�J����{���أ'#Eˢ/�@D�xX@���?�4�(�z\��u�h��\=]��|�Kɧ�zS%����k�ՏaR�F�-˂{���Ye�,�6�2�y̒�8�C4�&P	��{��ĬipBWx�s����?�֭;��_9P�*�����Ă��iNl��+��
s^��vmt��}�^��f��n=�TT��#����:�=���P�;�ݜ��y6�`��}g����k��T�����Q���R���h���	qy�'�}�� ��fV�`�+��̣Fs8�;��?.Q�p�`o`l���4�I�^��U�QSN���ۃ<��{��/ʾ�1M�}��橣�h�0ߣ`�2�x�:�9�<E���T����\wH%��R%~��m�Žԉ}��2��#Y�Mb�N%G�h8�bIH�`�$@5�,i��v39�(�c�$&��J�V��/������#�����7��c��J1S/R�$6��Qn,I�с��)�0-|�%. "���n��n�����zP��,yi�<�4��פ?��p�������@�Q�~a"�Z�u�er�3(���|�O��m���-����Q7j���,77?>�-V�������,/>Rs��1y:������*ۆ���M�S[�@�~.�V��K�xخ�IT6Z/��υ�e�H;�Ս��ٕ4乙u���<����Ob~�I���u����Q�_�����`�_S l�5W��y�f4W2���(��fmW�
�s��
k�m���̘�{��s���.��٫�־+�7�(h؍ !<�;�'�Q�%$�FÏ7 �0���o�7��zŏCQ�o�}�\����z���ԴJu>A@��r��V`B��K}�F��r�|`%��^B6k��y���o���i�Ǒ����۶V1�L���0*W^+�܅#�8�0rQ���\��I�����B��Y��8��2�4��K�mFI���'�<��&M)�T�L��'��"�+�d�pAe���{i��?���?^ܧPq<%ϖ��K/���cK���#�/	)}�ET��8ف��
$���z����jT
i�5�����?k�@\��}5���JN���K���'����F-V�f����pd�JB�� ����"�Y�YR�/�][M�b�w�j`2��$m2r�&=�b�$�n������ݗX�H���u�/M���oG��m��>�3�9�\�9�);��N�^�6�Ξ��+ SP䇜H��Z���s��V�`��b���~�"ۚ�\Q�Xi���wLV컪cc<k/���N��Fc��M¿�e-H�j	���8l�`L��g�W9mD�A�/��p�~�e(��Zz ���K�H�&��ä�Y���)��� lO�%��2`�Lwe��dI���#�`��?��Nה���<��\"���/��⡝���}ϥ���yV]�H��b��*���8��|�G��ˤ�hX��b舢p#VKNd�����[7�	"�Ue=�����0�3�}ִ�R &��z�`A��K͏k7�	rb˪]�# >�U�0�/:Q��jv[L�S�a^/��u��wwazef!�	A���"*֍Of(�^3O�f/w�=���{b������Ï���4��M+���-��&���ru3��w�m¡��+O�1>�>�k�c�r�uq�^R�Z�%�	��0~�	�8N�]bV*3�W
� ��� ��Yݞ�HA{�����W��"����ΠO�~��2%ii��ӏ�-�0�E��
��8kp�	��L���Ȅ.<a&�V�'��V�}a�l�e:�&��x���p�ɦ�ǎ}�ʚ"�?/�=��^6�C�B�����<՝�@ PĬY�sM��a�Z�j9�k�h��d=��n4a�GC -iϿ���.��n�|�!�i�|�Nf�nє�[��q�S���v�M~H��.�J�\%S� $pgy�u��H�C���T����a�B�a +.�S����s�w|�*��"���	-U͐S��HĤƤ�a��+�!~SR�ɴ[����%�T3_�E�TW�mT�A��T�矜�G�w?�UJ�Z��Ce�W'�l,}�T87����p�@Y��ţu���]_�A����_x��ƴ��w����΢���]x�g��7o,�#<2J�<�����XD˕��	��d�Cj,�TA +ʟ*�e�_0r+ƈ���E��3��,5 ��
y��N<+\��������Ӧ@���7����"�7~�m2U�qq�" ��W[б��_�D�8A��%P���z���5�� �_���x�L�}�y7$X^Q�p!oר�q��N�r��B�~�f�x�ĕ�O��jw>���T������c�c�vZq����T��?��N�j:��5:f
�hژF���$��Oj��^j5;>��/	f9Uz�r�ai���E�-8#	�MbC���o���;�5����Wm5c��(��c�["��;�Tb���C�9�%t(�`��iSU���X�{�$���;��sѕ�j�,;���cNH��޸��I���J<�X(����ê�6�>�%6������@�m)ߓ��3�<'Hޭ�I�5��GD���QKj��CZ�B5b�	(�ݼ��9.�ӣ�܄�~)�>�ȸb�^L&���D�Ђ���0����9:zFG�(U_��<�ӡ��1�pW>.ގ-�r�T?������ۻ�Nz�D4�0�=Ń��g�=2��bE�K�ϖd�2�횥���G�-V(�ٍ@iH\;�`1��en�V��i�f�nm���N�#�ď�~�_J���A��K=�%��Qd���3��┧����AW����>�Ƭ���Gu��P��[�E\�6)�x!U��0�b,�'^�֚��0�M���-�"e �K�-5@�:G��Ň����0�/���eYvϖ�$ {ؒ{(*�]@�SB�T@�LҕyɮV���]�Jl5n.��~Vj��=K�I �G�f����u�{���z��^ʰY��3n�Iuc�u��-�cN�c+ǍL�ҩ�`J��]�����9�G����'���G�����m��~(�jp�a�! m;�4�����A�g����9��i��5�p�_��*A����Jt��w�ǭ[��
�`���i����p�m���9�l����[2wN1&�:����V���/�Q�ͬI�ysi=b���$�L�2*jq�
v巌�}Ӧh��o@b��Oi���p]��@4Se��)f�w|Ƀ���7Gϛf��XT����qPV\���z���؆t���pS��I�s���Pe0��/�'"�7�x�[��=9g��r��n���X����"�XTz�@+��9�Ա&���~��_����t;�b_����]tQֵ������K���7�0�e&�K��7� ����G85���n-3��cl����?[GYؔ�=Y�h�$?9� I-�y�� �_Kb���5w:
7
�~髝�K |YJIғ�c�s���g��4I��E��-^_Ǯy�j��C�Z�8�呰ڴ@���[\t�{C����+Jm0��>c�8�6m��%�Z` �م�ه0_�������q;N��F5�cH?J)G�ߑ��׵������_��S_���ӄ�I9B�\��N)dZ�l.��Q�����>�X`D��)�
���CO@B�D�Ā���_ );����R?D�`�0L�2��y1�����a�e.
];7�!zHq&��i�ԆYH�^O��1s�!��I+oU�OUy�K����s�j�㠄c�h�� �x��pp�B}Q��4k8x��[�����]��|!,�>{�&��SW��i��U=e���@��I��V�����uTLNEZ�ﳾ@��J�NA�۸l���_�D�
�Y�RXؘ3y���Wq���#�19���e����ą/K%�<�༪J�"M|�����A�g���>�Af!>��&z_-d�h�̘@�M����QZ��B_5���oBQks�(Yb9�����+�0	b\#:��/��ӽ��4=�!�Y���%�s��X���ߴ`w��_vZj���Z9PV
&J�2��;�@��󸰖���_L�%H`��~R���H��������������j�*W%N&Ξ�ǝ��_�>�G���@��\Rf1Z�,ڶ>tIỈ�WA��2< ��o�*O�d��L��,�sw���F4j�z_Z'�@S/��	��_C����XdL��?؏*�p�y/F�v}�9|����k'c+L�@�a��p��YQp߫>���~�r��f��/F���=�^��
;�Af�3$�	�˾�aa�-a�vW�j[�U}�{`�xd��b�b�*�g�\=8^#����2���.3���?��i�GYό���{B��%�vȘ>��O�$�P´˻q�J{��x�Hf�;;��xV~��JPr�3h��6M�_�B�����g���\�k���0��(	�>	5���c�}���Z��t*�e�\���ΰ[<�,[����#��"ׯ���7߆��]�>AP	�<��*R�OϏ[Ml�@�@�MJ�����@�LK�p2��l���!��"�Ó��3V{b���5_��z��4>��������'�=M��
��[����'Ld6�+[$�����t[qV�e�2'��i�]xZ%^��ӄ���5����<!k�U��S����c�DT/�4�ڡ�)���Xcv­ϵ0w}����\dsv�1�饖�>��[ �_=��f�$��;���^9��]f��� #^�v�/k��/׾9*��w�6e�C ¶�Qõ4������ #mDo O�ˉ�� "ydh�ʝ#$<`�I��W�Rf�A�R��ϩ'-���ʸ���y<,�f��(tO����S]K��v 3�5�@����Y�d�@5���c��Gԗ=������bEj `�,����ݽS������W�d'a"�>�@iׁܶ8U���^)�l��澶��W)5���<r�:�ܺ�֣�4�X�'$�G��x?ҀǮr:tr�x��w0ޣj��?�F�0j��:��Qi�j͔8%��0�ԟؔE������煋����7F�l:��X�X��e7�P��~*xvJ���M����!�D3���e����"�
�i�vG��V>��YE��vi�(�Bw];�x$��z4�^H��X�7��ڌ������������4��m�Y7~=*���H����Ր���:Q,�N��z��}�XFQ�1�R�N�z�5kʚ�%�\p���7%'HQgnX'e&��(����W褢r�N�A��n�<���)��ʶ�%��F�����ot��2���1c�+�@�1����1�>��;W	;�D	,a�Έ�� Uw�15�_7�
[��br|�����1��b��:��kY�cb�V����O �Yh)���VM٭D�'(��YO�9�	N��3�#M��F1?� ��=9� ��H��,2���[�8��*��, g�-׹�����6����oi�F���,�"�(�4�E�[������vۿ4� �Fq8>~fwK��Sp�.�$�fN��G�l�����m�s>B:����+zD���`�2!� �]8���`�%l��sciG|v�0�9�����d,�	�G��ke&�w��b�x[ܔUT }e���<�ϗGa_������B~b�[�a?iu8]/W�ȩjS?Hi)����0	�?V�}�� �m���-K���(ԍ��`hl\i���[�}��C�h�����.���q�N;�����9�����`K��l�!�#��Ԅq��.#��Q���(�|�)�?���)ml�Y ;I���k1l���H��1�7�~�I9l�K�g��~Io]J���Z�[��k����&�\�e4.�t v�Ĥ���R=4��]jhw2&��<g�wb��]�5��|aګr�7�Ιv�a#gs����_�Q�AdƼ=����g:�`�컑���3���,����{`�ӫ]뾶�/z���.|̬f�����B@_�}�EfIZ��(/\/���̦|��3��3;�@T�=��P�,�Ȣa ��o{��z�@��!�f�l1(,�<����
PA�yU���iH��MU�u@k6�ի����+�i�b�����3?t�Ɋ�Y	��1�m�X=�-�n(.�`�^Vd�2<�5�(+O7���_-1أ�zhu��^0j -��o�"Ʀ�����M��:��s�5�l�7uˏ#�Wn�#�t)fG�u�~�K��@[{\n���y-���@!�;� f�<��r�K~J��=т�����%V�_��04���H�`Ǵ����gKT�K�(P�μ��T�/ܢ|ݻ�\�2��P��X6���2�����8'[p[����?;!Q�ΰ�C�oV<����ȠGUc�v��l�8_�;����ċ��R�Ĉ�����{�NE�r
W�[(���B�4)��_������N���א�.];�e�^�s�����yL0���i��z@*�Q�9lc*l)���5�y\h)0�HBv]B6� pud�1׎_1r��5������1�|	r'4�J}J��@�:��S��)]S����L��!�O���᧺ٻ���u�;� @��&*��>U�3.�
b(}:&SX^�^���k�%Ք/�uh�тb��y�{�2Ț|�ԍ��U- xR���}��>�s�k�����e�z���q!4ql.ހ���� '�����7���I�>�6���q�l��5"��~�qO�M#G���wL���h��KD ����ޤQ�\I��E�O�cVye{���K�$`qpm?$m�� ��V��%E�~Iڠ�|���P,?��o-$�/%����Lp�W��Re�Nn���z�P������ˆ��jc�Mt��⸒*G��%�??�*��P2�nA����$ ��+y��""�8��q�U#��h�@�G3G��2��M�a����*T �B��.g� h=o������pӣ�����3��J++�布ɡά;4�fı�'2�O��%�S�97+���ˣ��*���o���eRIN�*���2���Q�e+K�)�ɺ8^���c��us y��$��+��b���E��o涞��9:�����X��F�s#��R��J�3Yc߀	���eI��>ܑ"��=�x,����V� ^�$�@7��Aа�L,���۳ǐs��q�p�bt�/G�� ���xJq��J�XAf�#"�^�1����]�+�[<��C8h�HZ�X�6�}�R���J�>��ژ�	�7��Q��5
�Q�������P����\b+L���L�t3L�����9I����\�Jb�3�Ӳ�U����{!�G���p��"9�`	�¥'�+U�Sɉ���)�?PAo*ų����ź�[s.cO��������Mвij8J������"�i$	S���,���W�����M/N�����=����\���~�>�^(�_���GQ����V��k����ѕ�����=3*c�M��]�j4�uvPf�FzA溑�m!��~���~d��c�6���<���OL�A�����[^��W�3���	o.��[�a��#�sʆee�h(7�l�������#�g��gFF�7�"���/�y�~��ĬŜ�4Վ�lbQs���w`�Z]�Nv����Н�R\*]����z$ݙr�����ò���>������������ɴ��w��O"�5��LC�nүʀ�E���q�d�Ϣ��H^ 0�o`�D°G���X�� �f�q;�1u����}6r�K�3�M1����SمMX��'�m�g��|Fw�� )Ĕ��'����
Z��>���K^�ুP��p�8�H���_����>��)U�\�cr��
�i�3�M�`����W�}�4�:���!����rՓ<a��sj.g*�q=�}j	���=��\l��F�}o(�~��{	��lg�*{�&�� \��t��^��`���FC	ѝR�zP:�.A�X/�N)�(���ʹ�]��y1�{F���DnΈ<�^H�Y�o��y!��oX6�- �1����!��>ǹ�ԅCeS���"����h:(�H��f�
*�Q�K>_�s���D�ck6�"��w��+��@��&��ik��F�?���ae�Ak
_h��A�6;H���e�fT���Ohv�_�A�p��0e9�=gvk���%Di*���Iر�s-�6��w���)��ӌ�����᭱o���К�����?�a|?�K��WIK|��z��)�ogI�A�@6�|<S�u�djGi	�}M��\	-9�u��ĭ��.�}�k����MJ
K~��Y�[�[�����V����/��KnU~=.���	�+��;�s~m&({��I3Z�+]j ��BR&�%�5�a������S�n�+��wi@7�Q�����y�	�`W7�-�@���O�!����A!���Q�z�fM��T�S��?�a;iI��.��U�?�R[��z����(��:�
�[T��5#��f��Dt �F��*M9`�O�WJ7�q��B�x��%k��A���K\T[m�y��6�wL�V2��~���-U6��s�}�/�aB����$�Z �1�N�����(h��:�|D8�ӹ����L��L�>Y,�}y��*� ����c8�d���cΈ*[+������ʲ͗��ŒaR�-��;��^=��~��#���0�th�=t+Ckm4m��a�|u0��#�������X=��� ��X.���ְ�v�:�,���#��E��#ME_�45S2�-p�{f�W���t���\
[l$�V_} ����k��Q�Wiy�K.OV[���N��D�,�!{"�$ _ur�f�\Z�������)���a6w݇҃=�%�:<6t�ú�]��j��M/.�B����Y��7���jU����S�ޮ��#b�\b��,�b����둌`���6�j��)�������Jβ��H\��.N��oz)� _��-�	bF�t�z8�%��C1v廱�����S���:��4���K�G�~G��G�=$�7�#��c�M?�}��-��R�s�Ȗ���Ǧ�������9 �0�����*�c7�\��19��t�RA���n�K�#{��_�F�kwT�grQ�ӷRu0�jB�KS����0�<�q�$]3*э�A�@���LI�c���h�]:�숥[Dn���w�l�I-@�䰩=iH�H��!r������r�p]:۽*.�m�i�1�`Y�}(v"�pg<V���@�9��=�G���n&aaC�1�W4�� �;�eYC�F��Ć����NW>�2����;������J҉}{�5���Q#��<7�1��#��d[I���`���<ɺ���n�1�5ʠ�Q�"}t��i�i��ٔ6 _n���Zu��f�l*�c��=���r���=�fF�$b%�Qڣw='�'n�����*���L9FV���Cl8Ov�üȔP�>���co��;G �H�=U�W(�jDH�G9ҳҍ肭d�?����r���VG-��|��
D�}l��R%��R�;����kC�rK$��vZD��p���|��'샴�C0`u��+t�d9@�t4lS�0d���r��Ό�1��}2�3�l�c�u|�g�˩%C�FF�`u��΂K�>�}��6���K]z����)��zpU��� 
R�� �R���R`�[���	��#fs�3D���J�eL���*q�����`���S#��j�۽?�!�Ɔ���eJȩ����&�o�/[_�� ��i��}fB	��.�r=s��]S8�X���\+y+����� �>{~�>�߫7v)\���szֲ�v��0�}�m��S��_�j���u�⳥��a��:��1j����,x@�� �|�,�(�{N�)���8��ݧ��o1��
o����`ó_�� S��0��YgW��r��h��D~wƞ1"��.�-��]z��� ���t���#�4����y�_������z�����,>M���b�,�C=' �"ħ��t�Zv�¡K��7��km�ET�H�c�;�09J*��H�B��K�adƐ#��$�Zޚ����ul�D�LF��p��g�
٣�n���'���A8�j�p�S΄:b���*y�UU��r�0�	��s����M���~e����S:]��kf��o�g
�c�<�^��YA���f
��q0B��.�
H�������<��`�{���\n���j/�2/]��d�9IXё�L��-����7�U^܋��*�����p��uՉ�-)ʹ$�����dt�+Z"������6'�(��$N��u�d�����8������e�T�e�&vUf_wV!�/<�N-��,gX�>?Ը�<W��QGQF��0��>%��}Z- �����^��1K���zd4����t}��%JL8�ͭ����M:�`v���	Y3Y/�P�߰jze��s��X,��Z4���:E����&~�I�Mul����`R���w}�EɨxFj��V����1�]�K�� �ɡ]������EѽD��K7�c��������~$������f)�f/��jH�n���ES�}rܠ��J��عJ߼��C�k�]Ģ}�������S_��\7DIEˆ��[�YU�^�H�@�;My��Yb�wqSjd.-Sȱ/{F0)�l�Z��:Zy�`�H������;y��� 'nX���O|���d����W��<�S�� A�Z����D�<�
��uen�,XUZZ�g����ym���_��G��Z�:�[�&�Wh�8R��iG�;HO�ZȜ�i�|�IzD�T<�Ճ�o�������C�V�n(ou�Q������qe�PL�쳆Na�z�%d�)��;��4/ ���N|q�П��3#��}�����4GR"S������N�H�q����Doq�uC�ھq��"�m�f�˃�޿��
�kLQ�	�<#C���NfK�nC62,&���!b�7�&�7L��,QO��$9�*>����8���9a���#�#�-��H�����7�v-����{}k�׀����TL8�s*e��N`"�m��g�RL��v�F���_mB�Ky,��S�C�SbϪS������0����-��
�9���6�င�_R��'Tc����r��-v-b��F�����m/8Q��n�=\��C��.�!�4A���z�����%�
`�K��P��HAm�ȹ>^j�C�̵ N��Z&��YI�����Ǔ� ���-�4S��>��N'���+8�F{?�RW�?���غ��xUG��u�	�w'�X�-n?A �I��Ļ�����D}%�icX�;�����m��s�%Nؤ�Þ���s��4�谈t��F
y��hF���}�Ϋ��!���	/����vd"����TZ ��	*��v��B���+�Me����Aэ�$���+��%Ʃy��5�d��p��MKfy�����PZ
L}��`;M^D'�CL��y��$����f����%b^�S�����X��$�.M�����X��������c�U���L:yX��g���+AD�u�[�3a��	P+���c�!2�XmŶy�܄��<�|0R�m:�c�h�id�'���h�����$����;ѧ�I�Sk//�~�+#YH���&ΑQ'�����Y������o�M�k7R)�Y6��?O�m�aW���7O�5�<��8�؞��b�$_3zRFM�������E�j�d"N����z'6N��=�@Js�Q���H(�i���i�y~!�5:����Ɛm��U��hn����e��Q��&S�1mk�$0F~�{��:��d�c�)Á�U�C;�d>=��'�so%9e��I���1�MJO�ޚ.��㥖	n�]�/T�YNR���yu�f�������>Q�x��{���'�>ځ���:2�9D��z�I~$�/�>#������� 	�
D0YpT�k6T�N���$�o7�ȥ��g�鴛��V�o������4�}P��n$H;8�4n	l6fL�	�/I)[	iK9��|�7倡}6�8\EGb�(%�|�Z	^Ҹ9,~�9�]zIT�
��4!ؽO��.]ϛ��2a+Ī�.�l���Ѕ�;S�mE���:��_��6�6���t�8�W��v��l�R�\4J�)2���:��)ʤYΠ�������sT�n��L�H��;�r���"ū�3)�8����<%� 0,D3���VZ�4;yw�;=�t�5�I֟P��-��1Kx��<r���1���{I�����K{���~�9Wf1	/q�~!N��K[l>������c/�:�w7�!G+~��EiR�Ƈ�-ƪ5����������|r�]��l&1�^rg�ARwL���A�6�.W�8�h�\d�*E�)Pt21U7]O�yΧ�r	�����q�(ԓ8Ԛ�v��!k�]"����[N�9�lc�S�3���5G_J�p�*��T��;���
��٘��Dq��_2-|5�[��@o�idy�2�O>xi;5�4qwP/p\�éu�)H:]0�qcڤ�P�V��o^*������-ؚC6,�e�q#��-��sE�ya�0����I`+��SеPx~B^�����-����>)7�C�|$s�8��t��A�â8�!��]�͡�S(>�?������A"��ha������Y��.�y�y��<D�����u�<;�G=K�I�Qn��<.V���T��xz)c��j���i��EiDN��{�@�1MVj���ل�/(���9���H�L�q��x 6�X#�R� s��XKS#�%�o,/���e�e����ajo���C
7�~���
-p�aBm��D��3���Q���Ћ�-�S5At�Ys����d
Ry8R �`���
�w��,�t�	k$��m�N�'|���g�e�eU�G�� r9vZ�ً���0�@�O���������u�|��X�I����|!��bE���&��$��*���[�F(������}a?Ͻ����7zl�h��I�m?3&���Mq�������W����x��]�"դr~��������\�Ǘq�H�ti6�uq�Ү�d�.t~�{$%77�6��S�+��4�ٺ�MD r�f�����q��(8���N��҃g���-��K^�H3ۡ�jAB�c&s߻QfJ�KKv�8h
�h ��'���
X�L
Ǳ�#3L{L�shG��Ά��N�@��L�\�'#�O���z� �8q+j>�	��e�mD� ��i���R����g�0Xi�
 ���S]b��|�H�Q�� �?`}������Z|(V��̲�K[���/
>��%�����m��4d���k�-����03�V�<���4;��4�XkW'5i>�����ҡ`%���`/L�gF�0J�����7�+I�;�R`y�%��2w�']���?H}J/� *j��Ss��Qu ���Z9t(����헮�$a�U�C����n��`��-pٽ��~;�ΐ��Z�n�$+/�g�-�C�N��y�"�0s�n�����V����.,���e�fC[��@W�A�*��s�	1?���Mc��"��K4�m�yj�0�-�ew�����!��EFȼ�e�b�9��o�6a'd��䃒�I�SHW��l@��LS՚(o�K�3�n�x�%��ju���4�Ƿ��U�LŶ3��YE���c��5I=�3)k0B+��2'T9=V�R��
�C�mL�_�yZ�i'��GR�<�	HLM�=#�ᤠߓ��][ǭ�2�uȇ��kN^�7D��ė�̎�@��0�Z���cþ%])����6����|jH���.���NU���c&��e9k.)��T�n��c�B���3��\�iJjAe_+~Kv�	b����%�1<�N�]�PS5��o��(��� ;�}��U���g��#�%d|{��JQN�pGЃG�܊ڈ��z���.d�Dh�Y�u׼<<oى�Y�CT&j,�p�2 ���\Ii5z����M?ٹ)����)��u�8�@�P"�E��b�漻��]� �샬�Nd�����㟩�.� '5r�D�x����k^I)pmMg���L�Hځr�Z?�Z����y�?�x.��/���a���r����"ñTy(Q{'�!�K�ƻM2�\q縃%�5�7�N�N��ھ۠���CX��˯U�d�/;�����ckd�6�ٌ����������{6�d@(�� yk���]�6ّ,�16pt�
D@��������?�xm B $�ړ�h<<�S�M�|�`Rڿ�p��S�"Eګ�%ػ�PS��H�J=��_G�����|�ƐI�����L�4��,I,Q�u�����t=y�ӵ��m�,k�l͊�+	K"5���NA�}UD�'�0��\���,AR ��X]5 ��y4�Y`'	����D�M0 m�!��L��!�I���²�h"���^G?��j��¦J�م*�#�ds�m�|y��y�+_�&c���` �kn .�[�h��:EV�[6:��H6^uU	�4����&`��U�\9��;�4H[���d![�Y*��Dݠ�68M���s"ic�I9j��_���AL�J�Ӭ=�Z`�w\���� � B;m�oG �q� H"�6�yl��AM�1M���� ���$���v�OqO�+�9���.VB���H�x+�ӆx6��0���GF�!���&����� S(/��˃�����8��2���Ʃ�G 1"��6.j�+��K����<r���so�蒖 ��vf���
eߛ��~�{�j��7����yzmo����"��pw	�)e?�y���kA�.&���W�in%�G@�;��b�B85oa�F�C�kw?-r2 PF�^����OԭJ�e��⭇	|Dj|��g�z�2�&�n
��	�3 ���-��X��ܳ�,�.lt��@v��Ŧmjg/-�u�_nq��)�b�aR�m�|s�������K-FY��HSǮ�>sJP��*�0��zw�,>Lh%=�+�@�6W��Ysi'�?sn��T}&F;c�~ꣴ��(~ �Z�#�q/
�����!�t�d��"�Ri�'�[��͊8sLՖ��k�6'Rе��3_F�^'�ӀD���b�,��?����T)D`�y�J�ƌ��1�U�l�
x�'ɉ�f��KLg���6��2��r�u���
�����ﴺA���6 uЭ`��~bxTM��0:bv0K�IV�Zz��l�>]�f�`�K������s@�I+?Z���Ô���<)�[n��T�����4.���%�q+��6�f$L��������y;���%*ynka�i�h��t�!}|Kj�u<??b�B5��Xcsc��F�Ņ�|/�t�	��tjޘ\�'42"'�������g�X^ ަ�����#?m�#p�+�����-� �2Tu�g�$Aњhb7~�M_���>Q��Cy�9�u-���=C�?����mhlV�%(P/�$}���U�`5}w����z��b{�H�0W�YK���͏n|��A]�Ȁ�Ⱦ+)v{L���$��P"��@�?$'[A$;<�q��!֨�X�}��)��o��\nd�L\� ��8�@�v�	,�$ʎ�}�v�]JJ�hʸ����*~�ҋ�	4v���4�U����V����%�P�����	?D5\��^	Ӷ�
`�h���`�wQ���q?�I ��īR�Ч0�z�A�Q���ņ;�m�V�%�+�Q�
�����'�͓�s-��.�R�u��)���Ƙ:ޘ],sE�������o���q(C��xC���~�����1d�����0���D8r rp���#�q����˒���o�OKx7g`�E8_��@*4E7�E=?_d�!7x�{��������Wn����\��Ҧ��X��6�%T��ƃ�$2����E��<��E:�`Rס�t�;�.��'7л8i��愓�*'r�����ݦV�	Kq�~~��>�D�	)�DJ�o��/\2��|�-�h������FS���%{�e�	kaf[mvʡ�"i{J��1�ᐫ�=X�~���?�W�O���+N��J�@����-X���s-�:��i���-q�u���ڕ��	d�En��x7y�'�1z�%���Y)��ED�0u�a zK�J�Y~v�s�,@wCm�,w �}�N�6#��b]A������l1D�WH�NL@�>JqX�mB��� ��jS]�u芋���q�����T�Q�_�o.�0�6bX�d��z���
�O.�	*����!<U�Qo@ ��a8݆p��o��u	��pz7R��^ȭ��%�Սǋ�hvɓq�c$i�c�&���y�?�R
��Q�`��0a� mܗ��*&�7� fێ�?i{+j��z�������Ք�`�U_��2y��	� �.���]��5�8zc���8ǙP�q�!��X{�ֻ��}�녉] E�=P�B@�#q�/����� 2�y�y��ae��1T��н��y����:�p�T��iI���\y���؃�F�����!@	���iHz�AU5�Zi��\"�F��	Շ{�x&�,4�x�aI%8r��p�\�[�T����Ж?V��[hh��3�= ���TlԆUX\��Л>�|��^YV��������(&J��P0���5@�v�nC�?-�Zf�~�i�^��JK*�)���&��o^���6��&����~A�����l{�����h/��@6iV�I��瓶�#��4A�w�E��S��f�ɢm���C,��N��S.��0��W�'�_�4�yc!G���j�*��2�p|MԈ�I9-�\(���3��Z���� �+���D�O�@�����O�}�A�2j%�,Q&�D�a�::5?�[|h2K!b�}�W��]����-͔i��ׇ�{�NՉ�Z�~�����DU���}��WuH5�����pV��L�=�`J
����O�	!O�7��Ia����h��(Ej%�%�J�"����}���!5�t�|sU��.5��>^Y��,��8�<UnvhՅ��`�wb��h�ka�@��fZ�~�g��s�ؾ��I̠�ՌM���d	�Hsu�ה��ȅ�@a���|�w�+�9�~�C*"�P�q�j]o�ގ�qxy0����w�����8�����"���U�;NK�h��EP�Sxu�0;�Ya3�&���(���"�g��X�`�41D������SC=.ᮏ5၏���e}�ܦ��~����m���1���Xny���^6ј�~�\��'{EXL��8�lB]��}���t�����~o����X�%/��EfZ�+��]1�+���Ys!��¹��3��#�gT.��2�06���A=Q�㜬U~j��BЭLL�;�&OHpB�����>�����4ՠ���KE�J>�fց�t4�鴿;����]G�1�iŝ�Vj{�\�  'P��$̱<G�,��m6?�KS肽�&p���z��9��]+P��q�V�)�L��B��r�W'��f��%�<ܻ��8�轏�BJ� Gۀ�⪵����t^�Ɣ�?6�njk�Y�M��zٽ���E(Ş��X�]�)*{=��}�=(Vin��a��q0�e]������T%�������ѿ�ש����c��.hP��
A\o�����u�eZŝ0۽-^�*�9�$L��IxbU��9Y��IhGGĎ�2��c��$IǺ2�4�;�y/K��I�a�/̰�ꦫ8��"�Ӄ�������qG6��H,q�߉�u��TX38��;U ��/��.y�o�Ʊ�V�A гS}�͇��<��`�>*�[��U����7v�!�҃��}�f�*G
��{mN��x��-�,�����`j�"�F1�<!�UI��.��	�_���9�f(N�'iƪ��dg��K�@��j�o�A~�Ǖ���J��]���(�r�uP	WC��͜gL�;$1BvטG��}<w��h�n�a`2�`{D�W���Fwꆰ@Q�]l�}kU)�1�\ː1͛T)��
a$�:��oH&��4K�����Q򕔅g83�@��}�ܘ1Պ�2�c�*4��o��({�5�h�o��\R��M��ܡ��bo�Sl���H��u�:1�`ʇʹ_��,�_m�v�k��a��q/ɹoW�,l*��&˱7ezQ�c���3M��Ӯ�I��]��9��l�����i� A�J���L�_�����>h`hȧe���r\r�w/��]��OF���2��#�V|�=��zM��g.�H��w>�2���g냆������w��͎q�{qo�2m�,P�ʰ�&R�����A���S��c�af����AE�<��$�� ���[ZƟ@ ��,	��٧����"�o^��/J/AfQ�����tv�8�7P���u���]	��(!��oA�$�D��pE�7[~�v�>=-I��d&p���P�n��q^������
�94K~He�>kt���h�~xh��g�~Ԉ\F�WjIKH��(Z�zh��3���>�L��b�,0hȢ��壞;�M�����6��E`�}<{qU���H��2\B�*>�Z��[]�C�*��T�lx�ŞܒT���߰�	9J����B���K�����i�
U ����bt�)��3�KV��C�ȯuo�s5�����#�C�@&s�**�k��po	���B�Ac̉��Ù����~f���D��LC���g�伊_����Gh�a��.��OBZ��V7#�|E�>��ӧk��;�ޏ��y�ǡ��-�Ffm������1J�+Vw���6˱�ӵr��:|�e<�gH�+�9c<y�*�^|y}��;q�Q@�ӡ?^ݬoİ
#j��:��}q���V5Tun�y�kl�����E����k"T!zN5���u�'��A@8Z0o��o6M7�2�AW��ń��=���(�Z��?Q$~�Ui�G�'��n`}:.?�� �F6�(n�)��m���O�Fm����-�UrB|�0����搾$A������x�tc����ʔ"�WUb�LtZ�;�q!y�?���\\N5�
<�	�m��AFGU�{s$@�+/3T�zԏ<񭂏�7/o�7`1���XO�s��:7�˳�p	�P�&���#�/e{��ذ�	��1]t�អp�YB=^K2v���;��?�`�V;���$��O��G�o`7�a0���F��;J��o��A�#4RD�1ᢝ�����o�����tp��^�M�);WM)L�m��!j�D��ʌ��}ᶳDh�.Q���(�ٔ�n-������^
Ir2�r9o�L���#��G`4$�d�.c��h�ҋ���K�)21�6I�7$��<�b���n�,8�;ej4��H%��)��5�t�L{Ң�3�4�o%u�V(+��ZS�	�U��X5R�.rEW��8���~�3e+�`�."eڅLb��	�ұz��^
A���#�rt�e�;���\p5�"��v��\�Y�Gru~�6�Gm@Vfv�L�qr=bk֭p��QY�y)H�ԃ��(�4�'g*��ρ j�E܂����?يM��tM�d7aJO`ۘۙ!�F�J!��aRH�v\mO��G���`��*GNC�t�=�[�^w���EfR�.��*�q<�٣q^��JD3���&\NC���B���wv�\����q�ij���N��1塦vO.{RZ������P
?�S:����N`4�$EI3���ؼ��Ԃ����_���~p�ʩt&V��Bdl�{���ǒv<oX<��r��V$l?���$8���Kk��1{��d2%�������@e,�_�=�oB�_\B,���+�	*��P���n[>�Ʃ����8�j�*�PҀV,<�U8yG�.����g�t���>��w�k�C/��$}7��X=7�������+�}�e�]'��g���G��eVZ�������¢��壖=�7�LY���y��ѵ���sh�oe|S�K�>K@�e]���ڴ΄�-�ԊR�p'
Kb���5~�mBZ �x"��?���{��7�ԓ	b���h魗�)."��N��رZ�Cv�7*{ vFت����f;.�B�Ī��H呝Ƙh�!���$ɒ6!�#�̖�d��ō��i8�� cV��π{c�(/�vy������!������gt�œ��lY�dz�R�{�O�Ù�E�g��p�
��"pً�+n#�tS:e�W�F4b[/k������j�ާJ����x�:����E��x��5,�+mN��̔H4��1�d VY�Q���%�޸t���d\0��ܐ�:#]!����¶��6|�@��P���]����%��6�B��9�m``�ˈ����"��᝺͜r֡	h�;R/����KYkq�=U
<�m~#F^��!����6����T/d���DE�V��f�Ե'*�q`���sB�/��/����$o8�W���Fl����>S;�;�Oy���g���}2j3ZN5�a#���n��O*��� �ɍ�(`�`t�o� �b��]�QKP� �����a�k�J�m�E�wM�\t��4l��qhG��Érv8g�`so�\���I��)i�u<}M�~����ac�]�ͅ�i
J�rj�x'����L��`2��P��_�ꑼ{b����
h��Q�`��+������+�o�Y�0���bz5�)�0���q��쎽�"�W�4��"��&	�waO����:)��e�A�����c\�\�u�qH!��2�Kb#���>�TX���@�jc���k��j%&2�E��_Lb\�V[��xKb�	|��c�^3���y�Y��r���>��ո�����gj���x��� ����-��6������z�M�2P�H���ʿ�����1y�15����BV?��'͙��+^���c��D`�Ȩ��j�1���,�s�S��7x���׺�띧G*
�3�����P7��`e�!2�o��M�f�<�q����D&9=�����+IB��X[#L��'��T�hjM��q��M�k������?[:�����ֶ��(-���0\���⟛�*x\WT�j�S�	���� Ic=f.Uyד�D����%���\���ܖf}׉f�}�7���ֶ�Տ..@�����	\��@X�����S��NB|Y����2�%ȩX~��i�UtEO��L4R�����<}M�/P���'ҵ��������Z�*�5�B�f�q4ʉ�a�ڬ8E�=g-�������fz�(Ji�孊!�D�Q+6�g%�U(������6J9
�w��ػ����J���B�AA8�7*;�R8z���~�{��/~�X��)��mE���C�!N]	J��3��g����EJ��B�f�:	�mu=��;���o~�ly�l��G�� �f�)8��@Xj!m�9\�}^`�$L��Y�}"�U����{�Z�P��>�%�� -�GYd�|�W�Ȫ�u�ٚp:\��;�s��$�Y@��F��^V��#X�j�f�xdh��KS�k�z��~�4�7���9Y�*@�a	C���G8u�A�u��%i ��4A�G%Hm+&��:;�}W�]I!	�c�䡝�o�+��\�,�|�7F���v����!�������R�,\v7�vT���8=�A��@"ݦ@�v�mڢkr�@\7+F�Q5�lWC��;B�$�[H�`�$�PZ&E�ݲBJ�U�z����,��w0��U�M*�ڗ��/�}Ζ��#..0�in�0�	�wq�C���ב�j�f�'�ʜH(�<����*�?`�P��3/`GЍ�Z\cQ)���=���Q&�^�ϥ����� ��:T��Rn���*[P�|��U>��"ê�����VV���B͞d��� �z`#dڶ��*!�*s�_�P/�qT�v�x~�2V����ff���3��aD�S�PŌ��ϝ�,�4�GZ�mJ�������Jxy�SO+��t�g%�GE��帊A
&��1�"�k5άD\���\t�2�5�?���0��pE9O<�^�k�Rݤ�&�؁S����]f�����#�2�"��%���սlu���$wA����3�!�i���Q�R�r�D^bk��X�#����x��2	����RU���<@�֚5���xS^�v�']\?m�h
��5�I��΄�O�h��G�  ڃT��>dBތ6z(!��1����)��D��2�.wT,y�ϋ^`P_!�<��wRhz'�_�#�V���.�Z�x^��ƶ���w}�)�iM�'��H�m�a�ƴĮ��AT�=���R�-����;y\�#{�a��]�N� >pY���>�o��c����%��*��ɺ6�?�0�E�N�`v�p�T��l 7��:����i�|�'l?�	��������ǒH> Q�5�{My�-rS��qbUJ�*�y8�����}袹d˟�4�`�,N�>}f����*�z���a�F4����A{d����^����4�(��ەeƄ����L�D5�7E�th*�lR�ĥ=����F8��`�uT^%����ц�N��ZKW.�'�[[,X�t۫O�fk"��/<�����dvQ؏�g��t��=�0�����X��ǳW�A��l��*��j[���}.�i��	��+bw_*��j��s��vgQy�
0��o4#����ko��-l��Җ��?)�� ���ښ,+w�nW�p)QP���,�&
��G�R��YP̳�mGK��Gf1��	@y$�G��D�)��b�����M��3cÑ'�M``e����)����h�0���oE=Q���'6���)�WT�/�&�E3��e:Mb�����bX@��X����Y�G��$�e@/K�s���W���6f�Z#�;�:�4=f�pE��� �,(1���L��e�pm�_5Qv5Іw7��4/ߠ�� ����y_�uP:	���8f�M�!��F�h��;��d[K4.���.�'MD��լT�ړj���_�㳴
w��u�������+��T^�v�y�$1�OG�r�l�ۿ�KiT���f���C��y�_?���:�*l��m߯u\�d����Nq�нdt$���3*_��D�g�!�y�lB�U��UuU�믘�S��m�Z�U��,^�����;y7�)N���#�Q̽��kc!.L��,�ޮ	�=�^���k!��JЩ�_�c��;���^W�X�u�!i���׈#�Ir��	~;/A�[:�~����p?��a�ץ��2��[`s�-�����ƪ�����e����]���3�b}!�yyg}�2�\�_����d���n��@u�!*bt��zu�VXL����>w4C���� �
X��=������-�ƻ�&���BϽ����2H�������S%��󉑒\v�Ҟ\qL@k�� ^�1��	�x-�~���� :<��	uD��Q����I`:L{ �>_���i>���Փ�F���n�+�x��
��`B?���#+��]���K��z<����r̲3�WS]z��Z�N}�|��e��-!�DL9 fܲ�i�������Į�ji2�]!��i�!�g��7G�<���j+�����퍧�3�HW9\�5|�qM s=�t>��SҔ���s�?2�(��G�T"��BaH�y�����!2�[Xa�4f+y�N5K�4�E��i���~���5�	���7��7i�/�om��KT�����X�q�c����?��^Y��9g#30�J�,-��C��Q.X���0�ͭx���.�򀹬�Ԥ��z䇋%������h�m�������%<.���P�LU�%�.A!2� 8���͚����l���H֋r	�$��d.�O�f����o��s�^���|ŤF���y�M�%j=���ɨ�1 �G���5��㱣݂=���K�u�d�m�ܒ���;Ձ���ϩSP�v�+@�C~�!z<�^PH��wn���2Z�B�8@�<��6^��*
fM���,��ҧ��U24C�01���(���0���#��e�e�@��U>\ɽ�{�C�vZ`%.�A��|� !�ުwt��m�k�굱�mC�4�f}q�	D]u�T�za �p~I���O�����S|#Y;[<��݀S���׃�e7b=Q���x�_l/4���F�����{��g@?A<^=j#��0�#ͪ`��u�I_��
�^���'�� ���k�7��x��ad�t�Q���#j��[{��]�H��U��}_h� ޽�)'�������%�x���q��x^sKeCF/��&����񎝌C��u���T�+ŵ�ԛ
q�~}G�K %��HCQ ���RKY�J١1N6�u�sj0���m��IO����ھ�����_n�	�������7�}�;����u������Y�����Y�̏�xd1�͡,��;��I��<�X)�y�-��7���/&e��AӐ^ue��S��q��I[Qk\�M��0zct҆�����F�@����0.�nep$A�4D'�e(xQp=Z1!m�P)��y�=q���+L�y�*t�r��Wꉪ&����$��c�i/췧�h��Dܬ. >�p�/u�@2�Ӎy��r��H�e	�x|.���+oT0o_>9���h7�$ �1�N�FiZ��=W���3>���<č�5�0˫R��������{mX�8�Q>ċ{�\���"�7׻2K/�::�\QV	h��Y��}�w�������G�W��!�_
��]�����P(W�������a�$��NTB��8n�JX1��.��n��>Q\��h�s�#m�g�m%>#Ѥ�-c�Q��r�hU���-)��b�b��;��l�yc\����;�g�͎/�~��dVߍ�ж=�g=-�U�2X�L��)#��p;4����F��6��W�a]?�(��I�x��A2W/����6�%%��݃� H PO���3�J���IEP��3��aI��L��������v�q�2i�K�y������(1�R�U� ��"e�m����d��"��5p��;d��!
��hY�'f��*X��Q�X�߬���ey�D�q��k��		�yf(���}��L������bP��z�`nv�W��.�{'TE(	غN��F?�>���H�ȹu�P�#��������|�1��E���=(���x�:o��E��'q���o���B���Ճ��l!!|��Ģ6r�#�d��D'	�� �)a�`%0�����E��ڲ[��K��k�}�T�/��xw�
tR�ٕq���?t.�^�w��0�ҡt�~7��#ٛyδ�����Q�wҧ�b�����X~��Ζ�T���y�Q{�7�w{�^j*�:�mV��h�n������vdH{�%�e-�h��.�	����żIK��4��0�[ \<�����V5Է�\��Y@�+X��>�0�b�I��&�K������{�0�����?P�OD�P��
.����]$:K2�5M�6���7�l E�:^
��a�����`n�8�[1��a��0r6UV��ݸ͌ɞZ+�ق��ġëW��Û���ك�gh�y[V�:�Dk��tA�ߵ��(�
z`�e`���s&c�G�݈���jkʇ�����.�ڋh����с��ѣ�q�>�_o:ӽ$�Z���=ql.�My� �I4�_���m�C�������R��tC��j>���s���"�(�Ȗk!f0mxI�f�w4�t�Eo�m��23KΪv
q��m�Y;Mb�֠QT!уa���O���fr!���������%�	�D�v:�5�>�U��F:�}���:�K�/ԉbWY=,��K�3���UR�S����*�2��k\�o��h�M���IQ~�Z,�$M�ZFه�9c�t0��ˎ X�|�u��XH��oeB���2�k� �z�KY`�}A���B2�u�]Jl"����Ʉ����r{Rtq�b#��tfi�T��ł�Lҝ'�����BK����u�a(��?ˋӌ\���ۯy�����<Gc>�0��.)CV��V���,�:�g�W�����|~��j�?�慱 M�x瘚-�Bi*���>�N����v�\�27<��#zPY���X�-i}��
I���Urf�D�ʛ����X�'V�?|�)1 �.+����)`ޕ,� 3ͨ�
ͫP6n��7҉�$�n�7����$ɮ�a�{�T��!���x���`(ɛ8i�
�Z�e��[N���|���UST��Р :�V��z&lW㭟���f��oo�H���[��㓥tA��FLf+V�RO� �"��,�VA���~)�O��1����J�{a�;�g�@S%�+����|�D����Ȅǁ�c[�"�+��������)U~�\���p���g��⍎`R��B��&F��F.����ˎs;�����w�E'�d�>���|V���/���\0�ܺ	��.�H[~����g�uS�ƙj�3ۀ'�C�}W4����gV��i~�3����aV�$[4�7�x&��"�5e���Ƿ����m�jv�XU�@��+���d6�>c��gk�l�x+���%,A��!�[�
ʢ��K/���u��r�~v:�0���ݠ��Ŝ`U$��:��� ��
�6-FF��\�t����M'%+ti��g%�E�M9��X�h\Ԝj eʋP���[,3���S��rP�r��0�)G�����X3(G��)�^�����K
�1��43��ap4I-V�������&��X��f�/�A���$T��{�D+�^�X�wpd��ޭb���!�c!��cؓ�s�g
2�X������׵_s�66�e�^(j���(5o#f����sZ���չ�$�$��$x��Ň0ߋ�f�ge&��Ō)��;�K�^M�ca�%QY����O%k�w./�'~�
PMuҢ�-��Jp�#3cKJ�Hn,at�8W�Q���e�j��+��'q��t�l��()u�Zπz�����5!tnt,K���e�Ek�%�n;g�aH���Qɪ��W�3�"�����<�2$j̫6KbID�T�Hq��#�q56�:������A���,�[�6m���R/���	�"�=ݱQ���H`�fiҝqI�R��{����g ��|��ڥQӍx+��)z)�|47��S�q�v�l�G[���T�ʳle�l��i��("�1�2N�ǚ�EϞo�"�O�:����y	�J@<}
��n�<
�]�������]����ږO>J�|�]j�� ��s�#&{�����
?(oe��ɫCn
��Rd*��i{�mr�=�#��g>;X�5�	��t @Pig�2Ԑ���>;"+܏o�k�ʹ�w�yV�ȁp�J��h��0�_(�	���S��l�G<��-����Q)�Ҵp<[�͜2/��L�o���j~�=�c+����`�K�͑���kM.���6v�*Ľ�ϡ%�k�>�S����p�<�~�z�P�g�R�Ͳ�/��ŗj�e�8�z��\rݩ��39�2 �~+�^�Oc�� �<�1P~�쭝T ��pl�IZ�@�e��?ml�k�~ 3-9�Q��22��$؝,)K�������{L��È���-�!]����m3t�@�i��,:T��>��C��C��2\��8҇
���a�b�`���,������K�[�5,>Ғr�c�tiޯ_W��pL��;)}��c�R��v��">�2�����A�"��
��
�"���Eр�4l��k3�D���6|6A��9��;At�r&��o1�5��W�:�Xe��d�͍�$nlt��T|U���b�Q��-��8#��-��`�UP�mA��LBn9W��Ig���$k�X�W�G e�h��"�x�����_\Wf�޴�����B}-h�D�"�����Xs��7���G��L@r�T=>	s�Һ�Oմ���"�<�v��J�r2��Ʊ�'���1<�˶�����!:@�'�l��x6���0�KAH;!�`p��P�a7��iH�]�%�o�?��t8D�X {�6۴�x|V�w}X9R��Ԯ(15���;�2���a�u+`�@�L��qLX����(�(z��t�-�t���HAÁ&���c@gcƠ��oV3*Ғ+j�@�J%�$`�N�����4�e���\,LN�Xj���T��<l�Ͻ�,[�1 !������}�hP&v=��?i����]	U#�4#��g��D��Wy�j���􊵡kJ� Gý�pN�]�do�2����i�5	�wq����ę3�h��h���6�
�Ȭ����z2C>b�0ؚ�Qz �r=���q(�f�h�DZ&A0��G��i�.2���l8dIw�ra�-BK��>�G%��_%J�$�[�h�cN��M��<��|1R��,=,:5���@~�K�*w�4�d�4�ԗ����.��(�4�i�m������	)lE� SET��f����=E���|��/����#�F)�6�Ѱ�}5�-J]�� ���#�#e�Y�E,k��e�������yo(t��9T,uK���B󼦥)k���lZO���t�=�\]�}�
�T���^�i�����p��$-S��s�ST��C�Ul��O�;]�Y�,SRήG�v�3�2ZHX˻��hXiD|y��$��@"���֢W8�[R�}Y����#�2ٯ3js���(	�?9�턼���tjB�M�މܥY%�2z����HԻ��p�˵UG�Iz�a)V�C��f1 G^�F������3B���yζ�	�7�s�Z��(� r���m_ƣ��R�\�[�>z��a�� g.���7C�$��z��4hS��q���y+Ο؆�5���� ��b����`߶����	��4`Y6wB���3H[v;,Pw\fU���1echi�XsfTQi� "hN���� ���J� +F��>�TY�}��B��ֻG��U�C�>WB6	"a&���'���}f��J �'��E÷���Y�5P�9�p]�+6�c�c+3�G��B�^�S2l�H-�⭠OJc��g\6�~�/�w|kh�7
�"���E Y��K�
�G��~@5�٤"���N��p���xʦ�\Y�f&�G���c�zd��_��=֎LH�닍�N0��M���Ȱ%Y��C���c�2�&�~����2x���i�}\Х�yz>�0�����s�ʘ�b=aN6,I~?ӁG{�y�)�b�3K�Yd���t�Bn?��M�UN02�޵�λ�]Qg}]W�>0�6�k�|3�4�:�;�����IG��a��k�'�O�nOԛI��C�*��׃�N'������/��� �;i�G�e�Q-�џD��P��"Z%�k:����\wR)[}�K�C���s��3&R�L3����ϼ3w9�Ğ<�"^x��\���=� 8�Gv+�.0Β�&��!�7^5�=$�u��� -��6:�����(Rt�'��+�0�G�@�q5ziˉ�|��V1�?
Pc|��A�/�w�G��������TU�<-�Q���"��$PO�`Ż���|�F��!��Գ��4��X�r�Ϊ*Z\��%<�\,�k���dU���;g\�w��E����mH]#a�K���rl^�S3_�ud�e�i�RDқ�w���l�L:Fr7L��;��&!jD+Y�|��[�jGA�|H�R0��sd����wI674 e�U�E�n&.�b�N@nJ9*uJ3�?C$6��{&���s����F������	Y\d$��6@�<5�}q�u1�v[ѝ�y��P% �R�N�v@0�;8#O:p��8�o�5����L��M��*ǩh�$�6Y���z�,�%�X��7L�w�^5��o�ԣ9PN���<�<��K�0J�K�D���bv��3��K���|��S��^��~���� r�AL�/K��x�'�I6��O3?8�0$
U�HD���k���(?ނ�ϱ6��Į&�༽����S��$ڶ^�c����7�Tj�mZ� �Т�rcxɱ�딒/���D�YA�7O��Kn;iW�O���nr�'�'	v��L�9ʀ�ĝ�kqt"�>��N��MD�u��Cw:ҥt�_xU0�bL����4�L(SdxPW.9�;���~�/�T��Ҷ_�ҷ�ޢ/j��aŽN��P��x˕i,Mg8㱺�)�����Z�y�]9��.[�cQ��z�<s*Q���\����T����?���<��tW���Sw�s�|_k{
���<o�%"�ڥ��l�b�V�8��v�9 �����ΐ�ߺ���B�谉:5�y��m�,(+�>��1=\7;�	{�6��h�,N���l�4͈+��nZ�9+������א�nO�bFWA��$����3��Q
A��b8��*E��4}��d߂zBD(IM�;"��AA=#�IƦəJ�}KB�1,�K�2��i�dW�Ȃ����ѻz6��*OS�+�}�Ax�G8��)L�����z��kjR6�=��n(D#TIP40��nU��Eq3���.�I7���a�PI	���ݕ�&G�v��#ᗨ�S����oE69�{�9{[�⇽�D8M��{(~:z���]�j���6�U
d@W/̍�8^[��1���h�Z<�%�g�0O|l�G�r�}x��C���
�ġj��^H��.;X:9[z3�%����a�Hˢ�F���5��f�7��d۶���]�g��4p2���xa�����?AL�Ap {>�K�r"r����&vO�����s{B��Y�%�b4���&n���]5+N�V��� 
� ��Fٳh'�9���2�[�Y�1�����pDw�g5��x���U��cޜ�����m�����}�<�QV��;�	4&h���t"$G��}'�����AE�a/�s�Z�b�Q��L����I9��i%TQ� R�4�/ו1/ԸwHk�c�8*������HO�<M�S�=�5��ND1l�!�=��f��޾_`�����%`0i9p�n�s�q�@�r�����f:���AF`P�����]���Y���v7rcR#Ιk�¹�e�	ka�Dw�)H���u$f�?�T/irB`�R�� ��r��E0���<��������dƞpv�d�y�!�� ���k����;��L���0�Yx�XZ4(��}�b��x�7�#dN�c�0�`G�D:a��ҍ�_ۜ�e�m�������Kĸ".ʋ���d�84s�f%&X�Wx�g"r0���G��*���}į(a���q "Z�(e<ys���%��D�5�1i��|�q��D�ϗ����f�"B]���{�0��"���;\ҀB�q�,��˩�DRh������M;�ZU�㪻I?��Q�Bn��-���#��,)Y�]�X{�J���-�
�1�fz �
ܠ�W��?��!�pHPt�&���j�i6=��)]>-;Gt��w���ɂ$�\J$M��`z��4�R���Vf*��75]@��fJ���|K�?~٬��IkNO?���w���8c��;���0���WY,Y�ꏜm;��7bf��4Z��Lk�E���(ݨ>;��|R�Ҽp(U��\{�!�����T�8:��{�5�I�kH>z�*B&# L�`�ź
l���h����T�[\�5Yi�p�a-J_�sIL>���ԗu�);%I�����{�
`#�6FBK�衊xf�쐵�
��D�Z�X��}4��k/1�_'׺v���u��8e�X����]�αEg�x`B�hZ�y��������LPNJ�8��|m�}�BW�?�i��Y�EI�X����l�0�9W�ѕߖ�M^T�P	�	e��CCސ����N���r�Q(��ʏ��V�Tv[�e2@��V��D��
�o���؅�K��ǻ" Q����2�Yﭝq�|LcL\���J�U��c�s"��2?�nMԎ��nN���~�+j��qݿ�'�GT�n�J1�O7���.�C��)�f��u��}�<9��&�Df}-��ii�w��(�n|D�y�����n�	.��W;]j��>�H�9N���3Q�\�,%L[��u�u�i7ؔ��PQԅN�-c_݊�a��m��5��y��B�Rv��%yj�=cX^F����;��СD&y �h�v� �z ��ZK,ƉxW"IA���h���Z��!�	�]�*�����`[.e��:��c,����燑)*���c���o�I�¦
�����P���.`��}�
�r��8O�8"'����h#`�\���E�dx����nE���X6ID?�k�����%Pnz"�g�f�ǖ.U�Y��1ڡ� d;X�8�s���O
H����W���!�����`��17>hgָ4��H~>f�_ �7�IZF�S�Ҥ]~ި%u}����8q��T�Q�MI O���]-��#�n�f��	0w�Vm�ʗ[�B���_e{^
��ER��n}~��CE�<����`KY��db�)_?��=�I���q���ug����s���2���_���2�(W��X��n̤^1W�/'vo&7C2qJ㬢F������ݺ��C�D��$}U���#0���kq��5�"ߪ<2�	:�(/�K4+7j�n���;^ =q�@��,2�ӓe�h�C��ˡ�!���@�`m��W�V��1����D���_����C��G	+���֖�0}.d&�[b,����:�(8�~�[l�>��P[O���M\LL�h����ˆ7�\�E���EaT��=��'ٺ#` b����w�W2aJ�b��ݚ�� ߆�o�#�]/�Xp;	���o�&G��+,~Uq"�*/LX�R��[K"��2xe���H��@H@��L�v�T�F���Q�{և���v�y�N%{;��h�J��׫�+	�֤?[�F~q��}����0|B,?i�����]�X��KQ��)T��}gV�.b��T��\������RO�g�"  �QOGBėcYN�����u��V�6���	���� Z�W��s���:xԀ�կNp�F�xV�O���K�W��I,J�I���L�J�bq��h��A���X�	� ��:2-���e�]��h�}�ś�n@�G�,�r7"�f��rf=e>=q�2�Q���⺜6�1̯R6�ʛ1Z	n��w@���T#m_�_�FciN���{3�o����?��9�T�behGN+�_�R�G��:�x�-@ �9��U�-��΃7��<X��\���u��B}X$�u��,�c�A���NM	���n,�W(�n�g;�}8�O��f�O�m[r��n"����w���ʆ䇕�N���L�碿J�ц8 y��W��M�PB��_�MB���N��]-cΤ���`�$��\u_��cwT),�gV���	K~9�p�s}��	|��_�pz2 �7\�ҏ/pR���k(�WY��d:��~̆������`���-L�>|u�9*c�]�����S)�V��R:S�b�]�S(���%>A�izЁ|�VM�	F'�5��9A8���/xRO�؀��n�����0���}Ao�u��D�d�	�L���3mں���o��U]���{�[� �#�jE&&�y0[�V��K㰘�^f�|�v��*����N������?�YD�Xn��HpUh놓��M��]��:�����xw\0*y�?��n1<��aϯ�4h+�|S��'bp\�_Bm��掷���Ѕg���r�$n��>�: 4Ty�W`#��a�Wʩ��J���iĩ|�-�ζ�2�ʼ$� ����;b��Ā��E�#&j*��A�k9Xm�L�O�o�~C�񀸓�r�x�2�]L�7����)W�������1��bxӣ�_���ń��T�T!5�<�����'�e<�b��i��|��wޢ��b�TH��I���	�[dմ橒tí����p�x��Z�N&L��
��n��'�V��Ly|t�ek
��g랱-�D��g�t-�?��.�tQ)��K�T��׼�U������uא)W8MT�ZÙ(�����j�`?m�L-�?5��wśV�6xn ļ5d��Ry�{��f�'3�����~l�C�j�ep�\/	�e�Gm�^�m,�UZe&�R��77�p{��b�;��M��&���u7���'Fqb�1��9n�v~?\���B$X��>!W�i�����<�x�c��h.�^0�y9p-��|�s�dE���Yer�Mh�_����R�2<��jG��V���W��C�ǝ�ݧ�*"�<58X�E�ɥ����<�@KnaB����'I�7�H+{_��~/4�[�?�U��1W�nG�/�t����q�a4l��R��	�#�}PƮ�+Um	�z��d�?*P��z;e��G� ����������N�y���`����7ޡ�M���Q�P����\�AvF�`1	kI,@���y�Чk,� (PŔ�l���<0���E`{3�\5"F��̭W���0oz���[�5EVb:��Q6�8�H5�t R�hE��lB�Ӗ>@��0���0�����U�_�S��/V?�T��^��N7���"��pōb��svh�&{@�cǾr6xe�DɌ�]9�L��[�\Yz�8�]V���U^H"�=H�z�u��]���]T�����&��zf�|�pE���v1e+��Ɉ#��Un|lֽ֗�e�)"�-1�Q���u�`M\�h���'ʹ��=S����]|3�-�>�{^�C�C0M٫QC���A;�;R;�u��=*eQ(�h |���}H-v�-h�j�
��� (�|S-�Y��HSV߳JP���~"��:��O[6�p۟�v��������� {�=1H��奂�ѥ�No�g_Y&xwb��_��䭕�LB�7.� �,��	�O��U�}�D��5*�}P0�Z�k�v�d'A�����b ��,�;\���g��&�{�ޭ���w���5I���.g�"ͻAs���.e�g��+��m�˚Bp� w=F|5;�Ut�a�g�0�D�׭{�R��1�=ӵ\����<lh;��q<3���;v9��5r�a���Sקv�Hbﴆ#���:���?¿B�x����~��"�g�̈́+�S���]m3��M�^���>�ڱ#�����ӤU���W ���ީ�&s�,���V��E�?�˝Z�v��q<eA�r)��E��Q� ����v)��
�:�Ѧ��G����QY�VX�L6���31g�hf#K�`�1��U���h�ϩ���<���F�,0 �O�ő��{V1��rV�Վ����F<ߑ�y����G�u�w�
�H��o9�b�cZ���_u]Ύ�<���gAx�}�6�*Q�r�k� ƹx�ۀ �}j��5^���}9@�N+0�7k��d��0��ݸ%g
W	�
��'|i $݆c4����t�~q����7ԕ~6�������I%%��c��hq_o%&[�zÜRv��e����zC��F�v^�/%W�(k �l�YC��^|�gݗZ��;���ϡ����i��7���7۔Α�]K�Ir�H��q막D�	�F�V�d��)���?��}�_���%�~Xn�E}F^#n����j�lkb̘T4G���X�wU�S�pQ�C4�x@�tr�]�����2_�ITEd�ًh�ο0u��]� ���gԅ�o��{����y��Q��W�҅9Gj ��)��F�׫jw�:�9��Q��Q�9OcUe���;ӗ4Ű�]�]��c�}����b=)�OD�� &�T�ؿn=�iI�wꖭ�) �vA�؂��G���u����y.J�?�o[��E���Zl��S>��AnZq,�^��/g����wx;C�E���eo�vP�4	Ha������2/!ͩ���0���ٙ�7u����9���r疶>�liݐ��Y3
�@G��:�3P-�F�f���]�D��B�b��	~~�/��e@�꨽�;�?Q;�/�U�Ƴ���{��lS�ViZ�x�k\#b�M��z�߅��O����=���fQ�n,тo;�=إ;>U�/u�d��z�TB�����m��iE���[?��ܓhWUhw�JI��(WW�yY���l�T�)��I��r�㛷H���~�:/JHC��6�DVaS3,�t���DJ����3�T�p@�d&NNA�7�T�?��G��� =��؁e�Th�6�6�D���`:����g�fxټ�W��}�c�B�~��5����:?=��E�D�%f�7B_�/13 ���*��à�M�g'�7�T�1:�|�e�Ң�|�b������&t�ۋ��S�u;@��&�)�
��˂��w'Ě��Mr_�e�ޝ=?��Ճ�����̅z�!Ay�m�a_c.�d+���H�� �B9��_�
�eK�)��RS����i@��<�w��^�1W�Ŷ~ӯ¼���-��)��yd*p'��f�>��zW��6O�ݕ�ϝ��w~.��jl�!~�Wۄ@�)6~��B�c9���&X��[ǉ�� Ε�$F ��;/	7�2�#�*V�Ơ_!���s��s���h )L���H~k��;V2J�&�K}������K-���D��1���S	����~��>�����ے��$c����Ѡѹ����g����Oz�Y��o��5D�ǰ{��ۧ�80�}!�)Ps��"Ҝ��L2��!��+{~�/��p�Q�QB�EW�R��nc�A���`^��SIj�_�+e��q�*bH����ҁBY���g6��g ��a͚l7��q� D}�JDO	z#��6#�T�+^���s��Z�_�r��`$8��8��t�P�z5�3l�̅�T��%�LVY�`Dl�.���B(�p�쁇���d#]�5���#�}\ ]�a2� D�Kd�@�V�b
k��O݊���E9����K����p���W�/eB6$�6�r�Ed#���KZc�l���4=�-y�a�R���Kd�)\�ʞ넵�.�ّЋ< V����}��DP����}�m��0;9��a�#���8`%�فU�V�O��E=��*E�	-��ԗ)���05��l�`�ڸ�[bR�M�grg�m@�� 8Q,�v��|Y��.V�������*3�i��)�t�]��IP��z)/I�w�.��	)���@,���>����
�q�D|q𛻊,����}��<��+�� wc>���Ԓ[��4 �U@0gO突�﬜T��s�J�!ie�o���)����r2� ג֔W]��w�F^#!������pTMKO>sL�4�ޔfvf��7�8��,�Вa���l �J:Gg����G.�����v�0�k
���MbsKlP��JA�ƙ�zf;u�D�g?���O3~F��j>��Rޕx%�m@���x�~p�@y��s��tkǮ��M_��t�];c=�89�.3d��3�C�Ct`����*wz.Ƥu@[4k$�
���pa��5�����{%��'N���6��=��&HYeQ�W�̱$UW��&�$ފ�m����qb�* �Ǎ�^���S���k��a+u+���07��Ϗ��Kܟъ��S�ptU�DT��~ �y:S�nA�l�K]��vmXeͽ�e'ωf�\�̓����?̧a���
�S�����{*��x��	�v��T�>�AQ�'�h	yq��<�s�ȥ�o�(����m4y�zoG13��ɧJ|��J�^)�9��f����FZ�H��w��(�
D�7Aܼ��쭕�ú������|Y������6�#p�(ޘ^��]�L��>��6��Y��9�z��m9dCmWM�l�ra��'�(�����^g���]{�f
���t����B�f��lؖln�gB����m���b�n
���\�EL�f�IM/x�0b9�(�_�6w��J���dL�r� ȩH,0ޡ�Y�_�;�[��*�ǔm\�M��<XWg�ء�	$U7Uȴ����?��UUx�,����u�νҬ:��Ɣ��E	+��]�R�Da��[J5~�����?�X�EG�+Zy��(k5H�l@���'�̙OO���9��=�5��Ep�k"@K7ˋ��Iܖ�u�|��+�)�%"�o ���̍��!�*�k�캞�(99Q���$��Cr��c��2�|�a�bK�#��9h@K��YL:m�T���2�He�}�]��o��~����7���8���ĜI,�d����2���JMe�.$7��sZF>��K�4��s��ޖQ��D�o��n<�d�ّ���6;F;������@]��~���AO���[�x:h����N��G�ۺ����m �y	�#��(/�����Qw
la�|>S�7�}�1�Y3w�(z��?�ɵܑ�_lY*��u�1+��*��%�����f��c��iߚ˽E[�Z�dz-��jM�$>���O9���;'�8�[o�9����JV���X�%�4_�\:����Kes���g�M���m�7��x��7�%�&��po���~qs����}��4��ӏ�����{��ύLã��n�t��_q ��K���g�~Snؗ%$���/�S��w��9+�	�6��<Ѡ�*���อ��94��C�<2�>�����+��R�:/b,��]4^	������%<C����
��p��l�n�Q��ӏz��&�����fW�u^d2R?)�g荓 dPc���oܭ��t'����	�+ �-��Iҗs�7���SUY�8��%�up������4z>�%�̙�WS'�r�ʗ�N���GsN��@%��տ�SG����i2��c�R*��~[��D��jdW��J+l�"���&��<��t�r6i	��f��r��Jx�:U�J��k���h�r8�W��w�U��R�],�&��\��[���k��&��x6�~f��䯷�V��1>����p�Qx-�6U	qZX_
2�nnhyzV�e�/YqZx�Wy>�  ���p}�i���:�\��~�|��Z�u����b��8
S�V�XA��Ӝ�9���!I8vy��fˁ)�vD���G|����G����c�[����A��͖��������)�@�z�|/J��?9	��lZ�P�	C�8����̑��*I��Ί�<���c}yN�ռzhZ�!h19�"�� b�o��vj=ĉ�X�[A�8Va�&y�2�����y~X�%z����<�6/\��
֥�e�؄B%:��H��Co�?���%�3,
Yo0[(�����P~�m�j���m��޲�zg��z��LO<��Y�)�b���I4]CSJN��\S19GZr
������n�M�s��RE9����a��+�b������M�s��ս��f�[T�l ��Ry���{�����Ⱥ�1��樳dq���"𼯫!�8+����4�"Uc�*,��d����M��!��&`S18��,��Q�U��t�1����ٝ���7�!t�Ʌn,��+(KFU3��tP��ք'0���v�Œ�Ym�^nN��Vv��ذ0��L���ޢ�uQR��0�����m��ш#H%Ǩ�e.��S�ԣ���S�%�Zy����b���C�^���s�<�m��%t���h�]���[�[�٫�-}��D'��B��E�d]E�8M7��.�J���J����;�*�O����'\��}����Kp�?%���	����V���`qP �k!ey�X{�/��@��Z�-���P� \o�4!�{��z��'PT��\���u������F��!{̦�Y~�����{þ��]�fʣX�kJ|h���s�=��V	#�=�I��%zΦLr�z����vxGjA�Tq��|��~5����Y�|��yw��"�v��QB���0�I�L�Ù4~f3��%تD�B��px�G���#�<��O���%/kL�D h�-�)o�V��z��yLt��E�|���w�ґ� ��B�vy�G�0�fY���	Y�Bw.0��_�Bg�l8�����C�b����C׮�ZՏ��[+�!t���������'ˊ V϶K6�[[ka5��Þ�h��|}��?��2��[�����9ob�7�fpc���:�ݔ0G���P��JY��M�LJ���J�Y������3ܦ]
8�'=}_#����`��������A%me�g��h�e�>��C1"�U����P���`�W!r� T���i��f�weN	��I��?ڨ��{���&O�"���E}��V,�ܔ�:ć�Ɓ��N	�w��by��<���"��m����qU��@؝��y���um�6�9��g�K��M���`ߩ��7�b��;'�?L�f�E��fk�4�x^���k��wl�Qo���6f�8xm#ӷ�B�-������lpk� �B#��+=m�&�"�C=������3��#2�������s�5Ԋ���I�>L��n4ʩ�ݒY��e*C ��$��D�Z��m�N.�TW�He�V����u��.]�*5���,+K�Մ����
d�R2�Q'裦Z(⩤�-33,<�\�;�8ֻ��"����!� ����2{�������Y�{�4u.�(�+>L;ע�����1�F8P��yr1;,}/N���%��h3�9?�<h=�
^�ĄB&�����/d�5�DRL)O�P!6���EH�*�;���qf��m�/i���w�E���"�o_>,$�w0ge�)@�ג����חC{;Cʴ���ķ��ٸ�.�{<(S(kL�|؃v�k��m^{���ῇ�f��`�5�����s�)i�#�\�CyM�d�4U��k�>:����G��|na��3d�/"���Nõ_mf֜3�/џ�ܦR'�����)�d�H��jUQB�n�~�f��(�%z$\7��,|�WۧT��1��eRoP��hr�$l�����),�Y0��k�H�g�7�mr̹@�y-�E�Y��v
G�0̢V��'�()H��@˖n����}##�F�4EAZ)�	y�na�Ψ;㹟�����wn��ny��ndcчx�#�ޣBS%o�橦
N���Y����n�D|i���i�]��b�3s/���e�k՞-Us��Hp���/��b>n�����RZ��`�b�ᖀ|�D�,�k��hs�
Q3���f���W UcyV�����J���U.�o/�I��B9'�Y�ȸI�)����+�iG�Y���ܘ���%���o]�Dv�6-�b������4��,@�i)/[V�Ӛ
O榮�z���/\z��e0(� ###�.M�b	=�/��&lFzv�W�e�8e�":�rs2@a��d��K)���,T�j}z_(��J ��]r��7�p���R���l�@�\a3����������Q'k59?��O�u���Ż{p+�����;ȓE�t�N\�<NU�
��Kc+�y�T�'*�B�m���ߋ
�=��G��S��T�N�=+���EUQ�/V��U��E�|�U+�Sm�p�!�?�/ƹ����G�r+vJ�5��ͺ�^��#�Zk�����������&�x0a��̓�
�?DJ!`��z�A�@��4e2gu��I���!{'�=�b�(�l��S�\��y��Ģ�����.��l:���N�8&\���y��3���Z�-�؝	l�0GI󹝮[�/�=su�h�~
v�H�in!�bʂG����;P�e*���@KMx*PIc�d$u�}^�ٷ��r�h�˻T{y�B��}��Z��,��DYv�3���� �e8�=9���}K����V`'%yM���!Y6� �Ŵ�!cH_��i�����c��ԧ;�hq ��l�ape��[�;i�������5��ԯ��� *H�����N�)~��Rϓ��� pK?Q��Q�Z�K�r<�˒%`�`�S�L��/�`ڌ{�ON�<h��r����(j�*��G`d��f]��{�aB�3� �x��_|o$�c�#s[^<��0����]�'�
���;~%�`��q�>3I8�:+1�h���S��e��1y���f	�H��kmW�`�T��HJ��p��z�h�������§�s��N(B]2n�o��
�ɀ��A���jVF��m��|ꡐ�Jc��I2o��m�@:�ק��|�9):�39S�-��\�b���h,ʟ��������+XV�a��,��rȌ�88�'��c�ӱdpF*3>K=�KS�)�"�s/SZ�e�o�@`��Q���%�����E�W��R�M�����
<T	��ԅ��$Ӈg��� D{Θ~Fm�wK�F܎�h-"䛏���Ef�w{[�ͧ$�����u��oh�n����7���� /����~j��Ο�G���b����R����k��W?�J���p����V�:u�A�ܯ��4�:$O��������i�ص�>�v
%�J�[�"3���m`>"< A,�����0�=�1X���#�t���l�M��a�ap`�%�t�C{!�U�f^10�QRi����֍��#�͕����
,�uM�WI2c
���5#o!��͔N���ZM�clo����^��5o�������];\X`��`��a�
�����l+�3�*X�!���Jr�MW����s�յ} o\Vd���D�dۧyd5���l0���{>F��!���^�
�&���`+�զ�/��6�_��!�Q�9�%�@������Uc�5��J�mڅ�2VY@�H�y~�2G����$�Z����]m;F�d��b<����0����.�ɵ2�e�	���˿�8��7��[�H�]��}���KtR-^W0���I�1դ}�ĕ��q�e땈� �?�5_{��!���G�i�>���L|ně3��c�u?��&:�QP�a�R�a�9t�1��ƀ��\�����g�K_E��%e۝�������%�����T��4R{��t�q��v"[��8Uħb��⋃x�O��x3���H4t�����L
Sˢ���o/'Vo�v���v�|$rk0v�:a�
)��1�#Am�	�o�tA��c8�悒KE`�6|���A�����k	��9]0��H�*,��Μ�K�m��86]���U���7b�J�F��]��1Zd*�`��o�2}
�i�:D�]_,���ߥ�X��鹬91l,9낿2�M�4�V$}0���)��𧺵��)�Uuv�֯ ގ�G���S��l��X�m��F��w6�@,��Y�UUܽ�Rד���C���um=�q���wa=I�k��uP�{\��1�Q\��HĶ��&vV>��T1=;�In�u;54��R|�@�վ5�� �v�>e�ZpMc�Lc�
#Χ����6�+�p;�n���T�؝�����B�3=���\�M2���5d�Ԏ���j�O��������#����[�۬p����٩k�ge�	�������C��=>�`F��n �`��>�BOk2��c�n�����"HR�<1j�*-��m=dvFIG�x�J���I/��'b�WB{�>��ފ;T��c�Ah�i�	������1��҆�^V���x�3������+���)���PdNJK�ϘYfJ��|g�i��B�
h�nbI�s���M�o�ϡd]l�D�5=V�bn_��gGK��/g�����X�\1�Z��6�p�����]��a�~�a0��[[���B�c*X�Bxܙ�o��J!��;۪ �G�C���㧀Z\;�ܔ�v9���E�R��8�����Ys�%�i8�W R�#��vR���/�����`^q��� J��%�I)�1��ᬬN�������s L쯰 ��z�mD��|�
'd.��������rL�;�����~juzD���;V�
ռ���œ��J"�BD+%����m���^�xP��+�wJ�֩�$�"���-!)6��͙P����/�C��n�2ڳ���wݕ]�Vn�$��("T"�q�ow�r��;i=W����ک��){&[�W	r<é�x�$�g�� �z?�}�Kx���R�-H�j
��b��� z�����.W�� ������tXwJ
(��v��F�`1_KC0���^�*s�,�c9���i�<��?,<�"A���6��-�����\�m!�d���:Q?�jn'�6Ks��E ����s�C� z���i�R���]�[��P��������wt����k|�c�u��|�OX�t�)F�s����'�3�!�+��)IV���N�<}Mc�,�ЎŃ�B�o��uyt����Ԃ�'��H48��Q*�I���Ls;T^?^"����o��ʵ$1`��2]@s��!����K����z�駄�+�	dr�=-�-�`O\������0��+�� �@\�
��&|S��<�3=��kT��<�vo"���/D�`Ҫ�$�,��x�����#9Š���h�5����o����X���SϬ��.A��6n�%�,5�,���y�Un�&s�#ܦ�tj4�P2<ѕ�'�8��Ԧ���o��{r��r�FJ>���'��2o����v�!��ؾ�N!�o̶-�S[���`��Dm�<	(�|`�x�	�!?<�U��5�·"G3��Y'�g��˙8� }���f�p�@��o_қS&x͍\��vB.�R�H8��B�
�2R���XWGL�
#�
�4eSi͊6�jwAi�l8:b�cn��O�{c�bb=�C�i��G�	*C�1�yV4�����h�"T���	��9�Mv ;ݏpKB�8������6H��:;m%������L<�����'�h#���oD�8+$���z�	��O�!ݿ��ҊH�~���Cj�h�q�V:t2�n+�v�1n�q��Cp��v?��-t�ׯqG��Y*Œ�C��۱ t�ZԎf=�zC'5��̻�.�\�(�q��Kk�a��%y�:6T��uå����XI�~����<r���D=��4�p#ArT"ԃ��r'W�IlZ]1i�o9�<�|�S�VD)<��њs>�|��"4��i�}4[�	}����g]��D�X-q��e��7"8\7X�e��Kr���z��5J =cx,���uNe��a���^-��C�?��A����oI�u
r$nvP>T��_��ك��=u񐭘Pp�H�8�F\B36$��kR�9�ygB���Aj�@J��!��!�ES1��&��A<���q��\�6>U��Y�u��/�4���I�m���(�O����f�bPb��޵��&�/Y|�0$�׆GRQe��,���Q�V�.���C�E�����o;@y���Y���=�&`����|i�f��
G�	K�
������C#ǟ���9 [���h*�'��^���M*U�c�r|S�d��V�1��?����ߞ4�'Ͷv3�V�?��HX�?�"�����'\�.=�mi�_������[:Ah
���u?�u�)��'`��:O �hU�(f4՗M[H��_�Y�u_��G�(@f-V�sU���]X	�gVr�@����ϱ@�C��#V�w��-��}�>he;����d�w5��nH8��vհ�xP�齾�����o@c��3�E_�3cA(�Ef�����j��9π����l�D�)Uw��)5	��kG�zT��!� .��u�)���ff�3"C߫�#��E3�7�V�7��YҴ�1R��1#��Cd��]b�Bhl�S��~���w�v��Zz
*Q�y�ݲ�4}|��
sԪ#�vn6#vc�Q7,[�I{ڏ������o����mo���o9"d��-�4�e�������y���+�{=@����)���3�6��D�� ՠ�3��J���FI�F���#3e<vW	��[���s4�=Ū|�nwP�`H8!��r����M�v�4�o�e�Eɥ&5U20�AG�o�ssMQU��%A�Q�,F������QjΓ��)�E�Xܮ��_�R�:d�}ᨚ��M`�eZ�x]��]�����r���jH�u�O�ʬ��%�ƞ=TĈ�xzx0�R�Գ��)���?gc�$q�?��\
Mu�T�3�k�NO�, 9s�yhT��c�|73�F���~j��Id􎛷%+�gV�ǙRU7��9|N��s�P/1/�ܢ3��_
�\f�e�����oޝf�2k�LV��{`(�cbo{2��/e<�����;�o�����&�p�/ƫ����r�F2���T���K� t�m�#F��)@�5�]o��]7��&�$��Tymש&�����S�b�F��bώ���$-�}���b:ۏ���IP�p�}���P��s;kӨ��?*sknf��I'+�v�e�	tYfބ:���\.V�7O�I�������ໝ�x'�o��x��r�N1����)o(İw}��axL9[�Un<�c+�Le{m��ޔ\�:�����Nz�0ҵ=TS��ˮo��e�XO��=Tʦ5�6%\�] e#;�g�nP���a�t�Lb-�?�h!�d�tZ~�˵�����:��¦gh�37��p��Ϧ�B��UW�v��\�f�%���r�S]Kv��1�I��������*p����^\�#�1�F�=�\���Rj���!�p�"��#)�|%�w^<�3.����{�#Rlz<�������s�& /04
Yf�Ы�����C\R��.y��G��Ĳ_s��qN�*I01����|w�r_����W�� ��^�)e}���#{��u�m��%��5u��m���l �ΰ �?��n���X�!.|�A���{������
�
㙁�l%`��l���jT�QBDo�W�!���B&آA�Ȱ�	f6��6;'[a�����̧���?�f��Ų	Üψ��0����֞�wty�y3J�H��/�[�3�Z�GQ՗-��_���f�&AD�0���dN�p�F8���w](��\��<��[��_�:|Jp�!���=��U�̵���%F��
�X3_&�d�i��tg���D���)�y��X����<n��r`�o=��h�Vh��=AU:6�1q�|yzm����0w����}*"����ɿd|�� ^�r�__���V�|A�r]v-ļ늩	�[]��"b�
khF�D#۪a�{��� �f@w���!�{�@����R0�*�+�m��Qb��1�w�8�{�-�ԽG.�71m��]�2"N1R��=�7�_��B�^u���)��X�V�0�q7cy3�,�#��@=l݅s��#J�ʀ�Z"�I���9̼̘yS��-��Š��G�55�+�ʫYm�)h��EU���.�N�p�2��<B%������Р��p��9ŏ��݂7����Rx����-�`���力&ߨ�a�ei��y��1�|I�� �Il���Z^��\.z�U�N�:�m����@o�J��O���{�pTa*�G�V:-����T[�h��sx²�[��q��%��t�BOs�¤#?�2kg�Hd���[�9!@;Yanђz�m�����ܹ�'�H&���% ߒ�.N��lv1T�̇�P���^�dD����r�h�)韭��$<�Mz6��v�z��9���>u�m��k�>��W!E��ȧ>_'C�y1�Ϥ�V*������s�T�չ5^%"� g�GX�Ҽ�tUan��V-�
�ōf�/�jxo$��=�HRI߭Һ��zf��>ƧJ���A��#uE�N��:�̇z�����kX7��1�&����H��ga��,Z�;�Ӂ�t�sQ�>b������6�/ kt�������Q(�t��VONoZ�N<&f��\Dֱj�b���Jx����I�<����$��iP�����V9����B�-��"/��e���գ��l�q�|t�_L��|��m�ѿ�8�Y����%���/�ըs�kC�eIbg5�}!3��Xc�@j����b��>W&搳m<N��6'ǰ��%��[a�.�9�d���U��'oԧ	�0fQ��<Q�UQ���:��ܷ��G�����1]b�G'Uzg�5��ZRj S�l�^�F���SYJx~""cc}��l�p��'CpF����/���Y���1�Fv��E�����tإR�k�nE�y�p��J"�[NiO�����(%�$d����ݬQ2p�0�b.�"��m>�A@dB��va���31���ڗ��H��@�`�a��r��9z�>?(5L��t��e.�3`V(#ޣ(`%!bo�P�~��ñ3i�߷���S�À�PQ�2�BS]i��&��@�&PR��� ��������o8�fx�z$M����>(����-���y�)�ˊ���#���ZAW�O������Qrf�:=��.E�OW��3u���t/�X'�Y���4/�*�O�8��u��=����G,v����Ȓ�m�8�Yv۽
b��c�p��>,����{��(��R�L4�wy(���+6x�p	�,�����B�����g�Y�[�:VX��Ԕ��O�j����N�e_j�QT
V���kŊ!�&I������ރ��	���Tbj�S:�)�3�G~F���bf�7����L
��Ĳ5M#g���֔d^i�6g��ZY5'jG�}s(tAV�*_¾�~���`��e�F[[�B�P[��|%�t�֮\'�u�������2.�m��[=Tq�$��F)�L@��:�Ζ�@l��%�^�[Q��b�U�`5�/�B��k�S������I�;�A��
*p�'����:_a�&9��33�� ����IR�7�)3
\���<��g�mw?�p�FG7�E����X"˨亮əR��~�%]�U��
�\���CWj`��_�������I�j�{c�@�p���e��r�|��,�sQz��v4���CA�G��#��¡��cq��Ȟ}#�j1Oi���_A����F����Pi��T�%rE�`7�����7HJ�1��FZݠ����&�]`B�\�\����ﵧ��E�� ��_u6�V�ŕ�3{�r(l�9�kCe5�Y�d���|m�!��<�N&ăq�ս26�FT����+����(��Q��#�]��>�ޞ���5�I��"p�bf�vA��?��=d���&�a� ��*��]��{#�<G:�z�U���R��I��n�4�fD������\�~��������>Μ�۴��K)ֲ�p~�Q+2�𳂂L��e��i���y����e*YG����-�Ͱ�QqF�j�r��w6� {�	��y�e\����R�I���|z+3]`8�D�0���-��|6��X��kU9"~��DP<&;#aM~�`��tzk�VQCtow���`=�C��"�B��-@��k��}O��O�O��kt+@���lC�i9�*k�>�kD�uW)�-�Lf��O��3!�t3��`�3�8��zZ�� �?:��0�* Ӏ:��O�@��C9��o0�P{6����@��H:[�v�1lRV�T����:��2��U�kR-;0Z�/)��Z&\P�q��Y��^W��\���!����b���C���QC�d���������E�����]�C)��ɣY�h7^�2�%á��x$M�a^��O�|4�� ��l�h���)*_t��G0GG$ߺEE�3Ο���6*~��ٝ���It�Y&�Za+�`��_&�3���,�U�^n���x���K�"S5�D</�f��bP�#��_n��E=�Z�9c�3����\\�An��B&�C��h����O^������|FқX5|J`(ה�"���g��o���v�����gSϋ	��C 6u�k+M�h9���7���@
n�X��d�\�8��xHeW &,�:Gc�r���\�ƃ����[#�O��{���'�Q�3ɏ	pt)l���vx�v�M�pN���<��@��a�2��3۩-�u%��V��8OUD:@pl+j���vk�Xӫ�]�inS,{��n�л�l��D(��E0����`��=r'��V��(w6�t0m#.M[�,	w��[�'��@�0ۑU�Q��{f�����%��6�3J�jlo�h��0�7�3}���T��2QRN���S-\D�н/
�wMh�ħHP�u^6����턔+v��hbe� nqr /hȁd�+�kKX��'�n@�0�قT��B�ڄ�1~#�`�Pb|����b���+�բ��SĹ-���� ݈���v�LX�Yw-}^�i�Y>�|��bP#�n[dz�W��pr6��u�bi�U�����ӑj$Jڜ�U�ޚ�`9��")�Jf��@��&�n3ڋœ�t{�EJ���oԒ	K�錣��OpK���g\��e?����"Or�a�~a�9�Q�=�$� 䛞�2T�#���|����՛x�$
��N���K��;���UO@IuDx�	���0wV��$/�G,�!Nǻg�_�*��`{	�q�lI=�L[�š��F]A�,}���O�M94��u����K���]	��b./q��Lf�e���]�VF~3�F���� +xu��L�w�x�3k l���2����c� 2x�A:
꩷	��l���Q)����Y�^]Un���S-����Yq�uHf�����]�6��� �K8�����ZlH`����'WjC��Z`Z��;#3�")y|�.b	�����������!ʶ(W�s�4����`�L4ڦ9���%?P2�3�\�r'+f��qYE�B��
��e�9��$�<|�XdR��b�Q�xJ>�\#�-#)�/����	rҩ���/�$�cڼ"��ƚ��Ec��6֑P=}���y��K��/� �� �jAlH?��y
ޕ1ZόqQ�GT��Q
�"�e�5��y��@Q��>�~=�۰=(QhG��!�!\�^�Q�p�%aa$=��@�<
��%S(��#��m�C:wd x~�?Eזo�"�	�p��������CB 6I��,3G=5Q��@���I{5������}�Ը�O0.=d�;��-$p�F\��v�x��@��	.$J�`c�d��q�*K�<�T�5gY�_���l�d�^�6;L��Kڥ�jÖ�tRH,L%����?�،Ynut���Y�^��_m�+������S�A��K����+�R�m���l�t\!Ph��3�'�����>�|?����l���I��u�H	����J���+����������j��3'��y��3uSׇx԰\�R�+�6����iȏ@^�����Rv���3�6Ė:J�hl��������|��+N�����Y��:#����9ZcL�����4��c7�"�o���a�ح0§BY�Jk]�O�+[�|v�Aпu�S���i�Y��c��?����>�*����������#��z��b�vxcK�xо��爱aZ��#s��|5��t��Tu��5��ʘ��zY��g̡�],F���T�����r�OVd?��l6�w����R���ARAx;�����H2��OU
)�R���wG&ή3���"��` ������\�����x6ςh�H4U��5�%���k'�'�oe�r�YT䧳��KL�e�$(q���Gx��@�{��J��Y�_c<����l5��~��2�_^��X�A.��gŗ��3�)���O�q��=~6�8,Ϩ`p�g/��ӣ?�Kq��Ê#H4���|,��j����|����� ��fk�AFU�����:�9>)�!w��|�F�Hk�O1�f���b�Z��?��#�g4�7��K�lIU�9}||*�ǜz^ �]�=��%[u�H����|�7�\>�����!���;����E�yF�n29�T�;C�Qf�p�(LW�@�劳���K�p��!����հ����a�
$��:�X*�o�;<&�ce��1�ԃiɻ����6�}�F8xVL�d
���"��wu���a���lX�h]�{O����Uq2�U��,iU�w.'�~k�ۆ�p�ՠUZ�q��Ӕ��>�����e���M]O�W���~Q�x&1�-w	�a�P:��Ԛ�h�U��݁��?�]��]���K�/� Bd�B]������|��w{�_�U��-l������<�ä��  �J�>t��x�Y�!�����ً�)i��\��$e7��Wxdh���5yFk���Q��mԣ�A	�2`�����|�~4�hG���K���#\�]5�&'0u�V��)sP�q��T��c�P�H��	8�(e�ecX�������"8�\��X`��?�n\���Iġ�LU��@D
gg��gO���|8�~#���/ҽ=3u�HJh>���2�NI���9L���yo�̄k\�%�ٴ�3�uY/�.�s�JO�8̤��C��A�Я�_�G�PF�5#e���(�a�qc�ܲj	�kY'8L'T]]/��w��23z'^hXh[��US�F+�u?u<�3s���o�����hV{���=�x�TU�H���b��p̼����U�$bx�ֵ�P�kF�O҂��1$�����)���ҙM��B~���阌w����/�}J{3��"p�}�tx�w�!^�퉵��7
���c�
T�;���R �����t�hQ~��Sj?���dR�g�t�A���9�&��#�3�L�'�u97 b#�;�\�p����Dzx&J��w�e[�g�Λ[�B����O�*Yg�j�۵h�;��Ƨ�z����~oY���M��^�<F֑<��2X{�Hd2��F,}�+>��i����u��0� f?�B=문�qWb�i�4�p��	:�E��Kl��4��D|��iYp�@�W�|�4J���V�`(8vqSMw�d6��3���*�檇.�m��0Ë+D����_�Gu�ٷM�Drݳ;��㎑3d�.��L�|��y���5$�� T�qeoMI��x����� 8�k�kL 4�6�n���;����D��b�""N+,����%����� ��r�k|����*'Ж�\&��Cy��jf�P���e.���e���7�T�!��V�Ⓒ]����M� &�6�� �_ŵ��d.>�n:~^s���Ļ�	���Z��Q	���b�0�����δ馥�:��p=f����w�W��� ���u�F��tƝWe]m	QX~�HMc�!�M4D9�q��%�A{Y@�z����x�ehr��񚀑+IM�7O�q�l>��q��,h�-�Q�f�N�.��ALd��#���F�I䇷��ˉ��YD�k�\nWZp�H�}S���O�C�r�B!�͝W�O�f�1[��*��S�,���Olb˥�ۙ�z&��&�R�s�G������W����G��% D�jj_�:�&�0�Ơn�����)V)���B�C�Ěf�<M��ו����v�'e��=�i��L���o_c��^\T��)!I"�0�	�.��-�"���n��W�����+�bP���'���4��=| �VՐ�.�b�"�Qy�E��}��=�+�D�����:��F�6��Ifg�/������j./6�k/g��.�Lg@<����VpUr��ٴ��h��P�A��p3��_�S��V�&�_^l�`)��A#�e;y�����)��&�g�������6��l𞦳���I�n.N���˽���&�#ccXP5K��Qc��%F��o�vG�A���`��@�m�����,��Jk�<I��Iǆ�L����Y3NN1l���/;��ј��V	6bʐ�y.��_"�8�)���Nk�����G����x�k�}L6�Eޣ�A�m߈�$߆�f	�ů����rG�� %W/���� �S/ C�1{s������Lʡ�'�/��������B!Y%EG�sZjP2�j-���o?�H��V�d��ﾖ���l��Һ��$�a'���|֨a2Sd� d��WQ��)1�:}	�5���y?/�E	j/Ԅ�&����iB����Y�ľ������J�œiO��'I�t�lg��8�+8�����>��3��O�h�l�$g�f��y�j�����{�!������ϰ�%�é1�)f=iT�� 3�*4�\H�w"o錦}A�A�{o*b"��6~�t����(�`1�%ر���U>�0!J����L.ㅗ�����%�����3��Ӷh.{�ݧ,�'��/TM^�	Uwْq ��#F��6�-?{/e�0�]��OT1�
�ŧڧ�ւI(U3&���]���SUM;�w�4��a}�z��ڋ߆+s2T�c�y.@������}w���FD�ԺQ�� �pB_1ֈ�[� �kr��v1��;x����Qt��W~��}NE������Zy�o\�A��UJ!�[�Fy{��J��%ض�������P	�ÈY;RTu���� ��<�օl}a�d�L7Aߙ�N�X��ԹJde�rϽ�e �κ���Ju���Ed�ό6<�P?�z���u�=��C$�P����rM�Kq��a�!Z@^���aK�1M��F
L�%;%�>e�su�]��^pÄ�)��nK��2V��Ru͵>Qٲ�fH�kI��X��k�J��H�I���N�u��3ϻZ�NJ�R�T�Y�2���ܠJ+�E:ⲣa��kp-F$N��R��0y�t�{�5s��A���[c���FI��Y��hĭy�\����;�ܾ���J����J����8����n4���&3����xLY�XK�P�V�� 6�s�*��~y�0��eO�So�˃	�41���|�\38ObIuX	�����;}�i�۬���xs]�EG�Gۍ,� ���qML��r,�'D���'u���΁Fpq�/g=G�>�5Q_�O� �^�@����A��̲�}M�*�u{6��5�m�E��򚔶-R��*���^i�������1;��en(���~�N?���LP�"dM�FW�����)It�hk�x����s�{��Z����]��`#�ow����S�E@�>b�6�����x!�f#���G����!d�:dޥNTv��임<����I?�Dq8��7�$�U�o���Y��zQ�|�i�g���Fpt�"'M��)��ꎞ�Q��sP5�L�_U2wA��W�r��M�<�c�cDR��ّ
����w���o��MI�e�l���ތ��=��1��{Jsʧ�Sc��zϜ�l�F�,��T����*��`dU��~����u�&�?Hbɼ�-y��=@|o(��c��{٣F�-b<�����:F�AjE 
�*XR2��V�B�59����NK��� ���I3���ڗj�n$�/�.��m�e��h��}��<ZQ�?��@nu�F���)R��������H[ג�k9V��9��Ѷ�F�TN���c��4*M���F��R3�Y� a�b�hs��[�*D��\� �w�u�G�Ȯ��6݋v�Mִ�K�d!|4E^�~�7�^��O�A�	!�g7��'u���(ЖOaY)4����/�B��z Rq�ڭ��hN�EB��I�r�n��#��˴&u�U1��F��$��+ѓ#t�M.{���t��2���B���^ ���_.�Y���K�>T9��'��dˌ}�1U��X+������e}l�n�:R�.qS���g�B�<ѲF��o�=`s �BL0P:Յn�M��c�����P�jM�|ja?����N�0��P|��r�7�#Pƨ�=c^�E@�}G�n�20?l� 2�����S��n�n���E(��lLՊ�|p�0���a�ܚ�%�j<�)X%FK�)�{u]bT�՗�xX
ί�����%�u�Ś�@?>_��Db�����;.,м���y} �>�`\R�x��C���yMZ��䕂?�y���ge>�Ql�~�|�U�o�x��0��X�������MEb��O;4���	G3c�X=NJ2\��9�Y�xIE�P�`g׫	1w�:���{:'�Fц�A���G7~|��@�U2����տ����$+7 L�Rc�fĦ/o"�9[+tb�r˩��)R������%�ͶPKUa�թ~�F��d�T(aI�^VW�PJ�?�ǁ
"(���ռnGRȜ�x�.6�e�E-'Z h��&�\=��:��jkr�(U��K�%B��͑oS�ܫw
���rm|�i/�x�%�>lQ�0����"��(ctU_ �F��Ӗ��}fH�̉_RSM@G�N�;&B	N/-��]vq�b�Ȱ���!��=��4@.���Zܹ����}n�̈́t�v»�a���8�Q3PB���u��m�Om�V���r�ɋ�p����u�����r5�M�n6�G������')ot���Iā�n"�A<ćY�j��3�%>��y�/���G�0`�@揚4mf�5<� �;�P&n>ݑZ�A�1-7	�IF/zP�n�+2V�Mn����FB(����r���0pLԄ�������h��o����㨌�w҇¦�7�S�׎�ੴ�FpJ1���:���A4�+������P���յ;Iݱ�.;�@����1U��^�Y$��A� oT��a3��f%���V��M�]Oe#/~��ҥ�(Z�x��n"t�|b�7����o����qp�c��%��Ė���㧓�<���[v����y�:��? �g��4k GQ�"��nB���K*����H�h�b���Z�p�e�0p��W7��s};,C�F{cZ��9M8�Y��<-��+#hA<��d�(w��R��@������)BaDYP��F6"���9y�P֧#N�fϰ>�a�8�9�G}􄑩���	t��D���k��e(�R�r��`h�������<�d�P�	�1�Z܌�`�8��o�7Q�8�x����.��)h�Er�:]��</ׇ�L� b���h��'�(�[uԌqZ�5<�ڜ���>Yb""qG��"b������E�T��횚Z�I��N 9䘼��j��v�,�y�Ҥ�j��Q�NvK�m��ĿH��"V���78����#+ ����x�Չ��r��c�h,��&�vX��n��~o�"�J<���W^6T�w�ԇ��i��Dy�����(�ړ�l��c�'�ov��_2�,��p_*�=�o7.떲T�A�����}�{��!�	�0υx���z����-V����IE���Y�$߈�  ��e�K�/F9r�^w�ĸӓdI�d�w�|���"|\��C�;݅rC���E8)Y�kڔJ��<�j� ��1#!0т�C[Xґ`ޢ��u8�k�;�����%w�s_�NɉP��sh^��]�?�?٬\�mx̍h
9>og���3�:�a�z��YC+�T��n�H�l���(o��(��D�5�[ў��f��^�mQ$!ۈg��%�[9?�3gѫ���ӽ�F��,3F憳sb#U�r���A����ۖ��7V��u��A$�-��W��ȩ��:�l�T�|�bW�'җU�1�!a1��@���Dob��\->�o؝�zk���O�j��qf- ���FF
�])��Eea�UQ��C��Yݏ�.�L�1oߓ���O��O���.�
�͇��7�1���AG�o����D��9Ta.h��6k��^��-�~y(���}�ݴ�uS!�*��\)�mh'�\��?~ٺ��#Ze�z%;!�X�s�%J?)����z[�����12v�����8'>�r�,
1&n�K��e��R/�\�d�[�YoR&�"}u��@y2R��.x����FZ��B�r �e�P�^��ã�v���y�Pp����U��N�c%��ň�vb��3��,@��K�?,���op�>HH�\X�M��x�8��'sYuG���h�������2��h͡�`��q � a���=���큐�Is��_a��}��^�9�[�&�P>2�M��$-��2:���G�&`Z�^SƎ�l^�x ^̖+:uJ]O0��+pJ�􇙑R�6/�X�U>�R6_�l�J�c����A�Y���N9mȧ9�,Ē�q�����;NSf:���t��Gm+c���A�5T�g3p� ����[D)D�K�M�3F�O�|����mD(w���6�E�)7� 
S�&y2�" V�*lxYV�V���x���6x�I)�����R�J�M��׆��������"�����L?G0`�د�J\�$���n�]}������7&gC
���wu/R��c$Wj�ZfV���X-�Pr�dv�����H����C-z�QU�W���[�gO�]��jf=�3���
Aeڦ��Ra��~��=��^� ��𓷈��Z�"R��5^�ǳ����#�k'��B�*E~ ��rr�Mz�lLq�i��I�=j�Iv,��a�#V&1�C�N��Q������O��L�{l�&&W* T�3�� �}A�yE�(���4e�3���&1G���9�`ŧ����*K��_w��-�^~�U�	����a�CN��~��&������T��W�e�r�f�G�Oz�t��~����1����#�,�2SY_�4�D�ui�nZM/n���xK�A�N����C}���-��64�>���a�|%;�����!ax+ֿG�9�
ֿj���J�i��l{��r7m8���k6�|���%���M�B{������/�-���!�#|�aTA����%g��9^���+���&z���Q���)��Z�|N�O`ЄI^Yn��ot]-�x��B���-�}uR��#BC��h=.$��^bd� �@��ҎH�},�}�ѻ^h�Χ��-��P���g��S�v�EL~SZ��0�!E�o�N
W���D���g�.���¹6��eY�Fo�YtI���1�K~�V�׼���',l"�t�|z�ͮc�UO�}���Dj`,G����$j��ٓ�4� �FJ��-�vM����n�����iЋ� ���)�����y�#%I��^�1�m�mL6��PA���;3�'T����}�)��ɵ��Z�Ȏ�R�O"'����#e�3�sFe|	�֌���=#�YAo��Se������l���D�P���N1H�+ì��[���~�<|�
�8O�/�8�2Oo܍�� �v�R��?ۣ��/�W4W��K��3�M�6^\��`Sp/ud<u��B�r��Qv��Ǧ��"��?�.Rm�G�b|]��V�#��͏�����.?�^0�j�^���ak����X��ɂ،5�5�['��܈�`�ٝט���be��,�͆��p�]���D����f�(N�d�q��B���B�:��TI�����G�{V��7�RS��F=��Ad�͜� R�-�h�ݮ�K�����Z�y�ѧf���4=��v�j�К ���t[�hb�f�:QfA1�7��_���S�?�u|M�!�+�\5�Aq�O���׳�+����ܠ�m��������<h��&�	a�y2�-m��=���v�8C��j�G��ze��[�u?�Bഐ�t63�Z�L�i��g�����r�kS�^�i���Do�1lYȀ:�ez��]D�J6����c�l�ӄ����)�v�]?j: kA����˵�����u����������
N3�u�B�S\��,�.��J�
�O���İ{���/�<�.n1�|�M�X>j�	#�QBט�0�<�l_�ܺCIw���a.������kp�q���^ҵ.����d���i���z����V��j�\.�6ʖ�Ғ��2��(�Qc j\���I�ʤP�oNc��3�玹̦���Y>Y�Dvޞ���+�W������m�\�F���n
��kh|H����B��珬�pО�P���E(�<�q��di�m�-J[�TxP�� �f$!y[�awa��2��ҘC�/����q�l���[�Hd�F�
�K<��q,�#�ٖA#��WO�aj�}��ЃL�4�g�t;k���D¼y��N�����}�2�\�.��9���Þ��%�Ǳ��9{������� /ԏؙ>��5��B�'
͋���A�@0,5d��dl�򧺨���ö��/�Rxe�_lunj�qK}yMSu�ɇ=^�K��J�p
�j��eҌ0�-�o`�u|�v�z�f�M������d �x�t�R�홛S��+�ҋnu;�q7�D\�<�)���OZK.�a�v�����Y�o��XV-��a.������ �6�;&1����Ll�4�o�҄߮� e|t�}'["!ړ}���vN �:���oZRɤ�(�{n���:a�W��� yP[2h����L6�.���I/M��W%�{��4P�a>��2�)�����Y=���vb�,����<��qH�S���R�'}�P��(Pں
<�D��0p*�V�i������I�~�=���F����1W���=�^�͍W�{�]̨���,����Y��/]=����'�u��#y�M���ނU�1�p���XX1�
M�	��l�r�J�E��;���Jv�U#݊q�p%j��,{�6��i���{X�reS,cE섛��b��3n"8��}A��������>�(�;r�f��-xDXjC� R���p��r��q�P���g줜��1Vb�la_N�Ņ��AH}h\L� ��M��f�SZ� ��̇�ӣ��?�.�����!�M�p<��en^t��h 'V��^D��;�qn煮4�ܨ�兞�� ��]�LQZNV�B�{��N�+͂����751K<�&c&���sG\)^oy���k�t�?��ſ����zTad���sW�P^���؎7��%�U_4߹n!�!�VD�0��]��C�P��E�b�?��P1h�%����<
·5)g��k��YT��d���JE�d��G�D=�?���+~ӮO���~�2ۄ!c�:��&[~�e�=.�4�5��QCjD@T��d�/m�$e��2۾p�{<?r'�;l�M�I�����λ�s﫹Y����^aH�m� ��=i��tF��W�8�FAɸ��֕qu�E4t|��7	o�Y{2�E��-�݉�؁hb��)=�W�^�N�t]iZ�%J?��s��Z����hxL�jQP.\9?e֧��;���K!w��&�cg���My�Y�?��Q]�f7^�4��u/��?��΋�a]\���o�%h��&�L1ۥ+ L�����O���G9�+Y�J<��* ���7?cՑ�@�bԲW��\՝�(�����:Ǥb�����8�tv������O����������`�C�&stܼ�^-ZF�*{ D3����l��x��U��>����
U�?0�;��'���]f���yAYlΕ�8���l�A�����Ӈ\3�0�0ڂ��uDLI2qVZ��=��}>(&�(���BFf����_�ܴ]g�y��	Z��-\�=�ZVJd�J[�)-�iJ�#RLn34Ċ�SaY<qE�E
����S� ��tX
�]�F&�*20���
]NǛ|���y�M"`��6 E%k�@9"�{�r�H�XM,xC�U2k�g��c:۟"푆��=�pR{d6(!�pIVuP�=�.�+�;##o��/C׹���i�j�H�7�*J�k[�	rl�����@cli��DKW��
t1ڷ���v�H�};2Zr��>Zt#_u�ܘF��	�O���N�րr�ܤ/ж�+�z`��6�G2���Z��04csb0����+\˶W?��^�Q'{1��As;�X��'��	T_u������s���<#��Ǭ'&I��C�W�X���șVu?/�ֆ����{�'��û:�"y:���1i���/X뿄����
��79R��uQl�������ip��jm�?k��̣<>�+�P]�	�;��j�}2�
��7`��i_%��
3΀��q��\���If��7�润��Ӂ�
�tM.�5�%�A9s�3��Eo�g�і�n�66��2b�q��@<��|19A��݆�i�r㊎Y�A>`�tDOL�:`��27�$@>!b��zb�t�"9�������s�0���g�ȃ���~>�@-o]��fK��G�=y����Qn�ļ��-P���,����$�ˬ�< �S�\�dK�	�J���Sxgƅ8��}���|9���f	9����J?+q�R��Q�l-P�d��z����#-G
����;x�0&�K�<�<퍵>��}���A��۬�Um��C.�o���Β7�YM���g�O�Xh��W0{�����A�M~�U�S�O;�����b�>NwY^���W����W�1�6u� Z��\~�v�}�Ü�s���^$���q�eem�)��B���tb�MS_�,��d��:�v��t��iq>S<��WfGL�-��1%c�7v1��fտ��=V?���x� ���3�R`�k,�,`���6�C���.bz�0$߆��E�N��hZ���{��տl ��;��8����Mժw������s �T7Т�5!�:������<��J�������M`��Iv����u8u"��CuȤ=ҍ�6��kۮ���h���"�x`��$��6q<~�9�N��r�$*�~�s#�XlM�y�.N�V��T�KKh�b���L�������B��s�b�˦��侜���)��ի�ш]�������j����?t�3=P��p�9<���+LX�hŚ��g���x�p�egs���~n�{�o�}
�2{�?8H�<�~{��ee��i7t��Q�^��z����!�%�V�v�`����K%���s	8{p�`��d˕��R�\�8Y��Y�M�f�C��N*ps�R�ᒙZ�V��\�O%���jSCK�^�|�+]��m��hs����?ǥ������߉�]S3iyb�^�!v=#�"j�/�GU3�Aӳr� w������B/� Q����-:����Y&n�T|o'
*��)`J��C�y�I��L�Œb,z�Q��s�G2�ɾ�K����5�3w�3:� ��qn��:ܗO7���g\��M��d����d/+Sc�N?�}b*�^�����m�CyC���s��JF����H��?���'}	�o��Ƣ��8b[�pRZ��]Kb��]�T|X
�ҺְSc��.��Lh�*@�����n�;�8���P��'4�Ɛt� \(F�1����^��B=�I��c�)�*������U:u=��/��� C{r�|��{�*�ˡ%F�n����ԣ�TʖJk���@�u�Z�ZC���rJ�W	aO�uK��E�X]��<�+�q�+���&�V0�|2�M���no���p
OT|B�1�N�[}5ܪ��;t���R�Rr���ϳ�8
���`̗<�箯1���MV�B;���Iih͟���S��'N+1-�5ț��Ehqx/-c��J�[�[XV|f#���C�v���pǌ�;�gFi.���iS���DFa!�"�=,V�+q�b����:��w#N'@�F��P���l��� 
�;���T�s7�?lAQd�)����͟�/"+%"&��Tq�)��t�(l~�K�Z�r��6T
{)��VbeF��;h�p�.G+�	�MG~�K�U�6�}����a�P��^����ț_��s��a���ܽvC6��z�Vk�n����3�ԫ������B�ڤ@��a�x��2SmM��4nU���"	��+H7���s aO�%H��U�/,�8QJ�cW�'ks�!ܛ#\�M�U���)Ӝ`������o@>rOj���X�h�L��oU�Y�u�NTh/�u�Xl\S@�k��Z���m>����?�jZ�)����0�1�7�a�YSV�]��C �l���w`�pi�e���&�a�� IN�衪��=Wv����ƻN$°�r�������J���U9�����q�q��V����
��Pkz��n�%���"
jbV�Ʌ �.)�����,LԴH���Q:�.a�`Z�AG ��{VS;�;��eS�GgF��R#�2���m�j�����:��ݏ��j�g%f/RHy���ݢ<����6����g�&�p�Wbok�o�-���cC���q��"�.��T7�@Yn�z,��*{V�#�:#S���t�p'-m���r094(�6�)�,�;��#�$�K������LOe<��X�My�����7*~�}����;�1��+ˁ:=��Qe�k�0@�vӷ(p��KZ���� �GKڊ`aW�;��L�PRw9|Q��Фe��v-�勇�cda�x
�xv����bv�2��z�dy��<U�tGx�<��C�Lҵ�	��g���?��mnZ>l;_V�ِK���.����΅p`��نlY-ܟ2�+/l�*�)#|"���V�#�������ڌ�������¹` l�������>���y=���s�l��\����i/�I8���1�v��03)�ӪtS���[C�&^Y����h����j�]պGD�I���	�4	�Ɵ��1t��nv!�#o�{o<T��-؟�q����-�R�θD��N	�A�~�<ii�#�P%��H�u;���֙��u�n�I�g�$��v�G��[��9�B��&m�l�B� 1�� �5��OV^��#�:������2Ui�'�(55�]^��u?����P�<��Y߀!x���%�%�>��r�����>�|�Pj�lx07<�k ����Y�]��,��c�w%:&�!��e��^�\*5Lf���5���NP�"�t�U�<����k%X�Ҍ��Q�R��{]|��y���ʜ`���0j��Kg��q����G)�d&,%+
����4|����2�]E�C��9�n\2��n=\����p$Ym��߯S�����$). x(�ڥP_6���U�z����g��T@b��L��l�w筪k�Y�>��:������13���=.FG,RC��&�������I����S?��h�s�%/O�F�!I.-FH�b)�[I~��ʗ��`"�&����-�(�b�1X..�a;�L�s�7E��Hg`
���Fd�2&V�rp�<�M+=��ɮo���d�����|&A��:>��xG
���f��uć~�oh�����1��w5J���	9�yL��\z�	�;"fi�A8(}�2�9]d���>}h�rp�.؁�/@��<vp����Z���֭!d�R�U�NՉ��[�����]&�|O(�Ȑ-��)�	k늠.Sm�.1�R�Z!�5���E�Ѣ5R��Q��K���Y��^���r�V�ECR���؋"{>L��ښ�pZ>[�w�0�����K�<�|,���\tr?��a��G� �˼�
g�p�H�f)���nX3@�=F����C�]�>��2v����##u(��aV%ظ�P��"@�[0-��C��MJL����K�@�h�݃�L�%u� "��(&W9搚o��1>E`�fuH��Kd=���f D�����>JY�j��p�E�WUϪ0g��;��Y���ƣEdx��Hɹ��e�_�H�R�5�N���L�uDS��kP�e�#wըҨ 4�F�K-p@�Bf/Ԥ��р�]_�� �Ȏ9Q��rR�1�궘	�,3�jhu��ӯG�i�S)�	{5��Dy��х�BVĖ2�#�XB�B���7���^Bܨ�����\wx~�8�N�3ЊG�?�ĪC�*� _�b��4T޾�}a�o�����g��˖���\=7f�r��4f�����"��OТ����^z���\ i	�m����K�C�K`.�)�&W���]m�A}�0zE��Y��;�����pj�L^ʠ�괰��GG�Ȋ���<RqS���=Z��]����, ���1�~��g��E�ڦ ��`�3u�)uR����C�o!��"px��`&[9N%��j��Y��H��ӯ��za�X��'�գC�-����NH(8d������*״&�O��2v���g,�$��U<t[�9!�]w�my�}M@��T�^ �����΍����G�3�j�Vatn�))]fCZ`F�%�j�g�� c�C�T��fv,'{�3?�gx���K/�.W�,�Fuˢ#ׁ�?����a$(4�B.N-�A_G����Q����;���!�t�z��O������
���a ���IR�f�=��2ɩ,�]]͝�^���pΣw��ۺ�ۢ���<���Lp��>���&�1&�f����'��O�OL; Z˾N�sU��r����6o�k]0�B����S��p��ڮ��A0ј�����7��G��z��-����S�Z�V��^�����k���d���8�|�a�c	����Ԟ�b��r�3��V
�0*(�cj�4��%�h��9n���N��C���[al��ę��p�[�Ա���'�����s����6Q5��OR�y�E�k�s�ϡI�w�;X�˩�6���y��RPY8��3�x�,����P��N&���h_"X�<Gt[��S������$C�KmI��a��mЭ����vÂs������Y1�˶��˲���sqD-Y��E/��mx���t���tR��T���A���^Fv��z�b�ON�����<_�m�6�r����6�vnQ�g4E$�d�S�R��m�?�YEV�)���*.I�ˢ	�á��gۡ�0����s������rd�����q���D��qU�)m�
����>��C�+G�?�У)���aFm5/"G�b�i�LC�{Z�%�����kԹ1	Xw��k��U��u}���ٔ�;�Uf�b�j@�Q�5H�Y!����q%�n��~�?Q�"n�%��NQOp��a0�?�i"�L��B3\��_�,�&�[��v#���w�����D�>{�VL�(��-墏%9�X��b�-ՂQl|��Ӧ�#eȳڤ��ai��Wc��l�$\<���q]N{�T�'�tE�����j$p�3fb���@-��F!u57�[X%���0��;��֓`��n���������g:[��f�L�B�U���3r��wP*nIy~�O>��ߨ���X��ϫU��H�W�y�����g(�|Ss��C��9s�h�ua�����ݎ��U�/	���:�^���	�����7N���1���u�U@�߃�̸����Cu��"��\%۴��\�JCn)����3..����D��@�@~5��i�Wm��jF����7|�-����s$4�tKϿ�RH��Y����=f�ŉ�
�̼�Z���HZ,4?�s���=�I$�;�;�8=Q@����do�SF��Z��z�H���.��ק�ee�(�dm�J�p�hA��2���b�G�"�2��ߗ.�<��R�*�Tbj�p�N�����'�#i�?��7t�f��7�����D1�u.��Ow��*��t,c�]���u���WJ��m�A��k
>�Nڌ��O�l]�����n8j���L�(dΌii_6a������hA���<�]q`p��ޭ�W���>T����[�l��z�x~Թ�A�N�>�g���Mx�P-qB噞ڟ:�y�g����`Ym���-�6a6�q�iY�кz8s������(̗}�&x��۽��֚��
��v �	�/��Kx�lXNe�<�`r{^��W�v��������y�#uX��1M��Vx":�|�_e94~��n^a�R�Oo2R=��2�	n�6��,���\�z4�	�H07���Aa9�x�b�
����(l�J��Q��?_�N-��b6h�Ш�x���:�˦[.��L�^�d0�HS�]�����b{�3m�b�c :	
N������;ۺ��/�������)/dd�3f���߷�S�k�	��;�d�P�Р�y�4��o�ⓟD�ʍ�̣=i�y���eэ
	��(�[ ��t�jO+�;�`�a��ʥ,e��Fv#^���wN�ٸ��8$cY�+��A�+�P�x5�@_�g.���V��̼�2
ZGY� ���N)����E��1lX1/B�����u�C�|�����? ����5����vW����W7��c4N�y;ѡEw
�o+3�$n8vb�D��u'�n��e,�E�<��	�85�m})~���,E�-�y$ms�٢/�dQ��K�R�	yz��t	<e��*�í|����O-����
rtk_��|��a�0�c�<3P)��6�+f��-�j��'����&n���&��<���yh����:�w^1������)��S]��XTL�I��]$���y/wy����oJ*w��1��E�_��Vm=k=����_�V�	̳�3�¤�ev�O搄U���M4۴zU|:�S�w�B�͚�Mw��C�{B ��yFn:�^'�֤���9<�hk�2�����͏8�=W�,�A���:��CK(��� ��A�Txw/�D|/-�=�ⷽ�D��>��}EХZ�UÅ��H���q�]��_�[H�6K�T�%�ԓP�
��R��"`ۮ#a��W��m�g����Ջ���9e=K��O���aQ�����C����	ҏ3�����������.<��k,���h��'T�ZPx6�2�˄]O9�n3"O��f0���Y�@��U���h!�4�dn.�`=s֑���xQ�9���J>.��A�5��?U1N.�
,"z��D��~�U�*��N����a&EC!DB�:)�D����G���H�P�^��8���"�lG�Zy�P�3EW,�R��pn�|�q�.8�p�[px^ߍI���"�)�.���&�-�_j�H�sv����Wu��Q圶��X)�?�};'��3��%�zc���%�n��5�t����C��5u(�Lڎw��](�d#Y��V�N�)D#�Җ��/�Z?�����`6�"�I�Zxlca�ږ�r��NG\�t�HL���.�+֚��=Ѫ����|�-��5��PO��T����:?<DA�ꊷ 05V���=���,��*z^<b��-�0o�F4/fi� �M	���yJڇ7�*�i`	��߫�Q(*@}޷Ȝb1.��%�<�c�i��-�8^�$��IzYUh����]����rVY���>,��M��Uq�Lu
��R�G%*��[�c��*UDV%�ăH�}]F�1dR� ��q�v�������`5���P������F���r����.�|\�����A9}	�u0��X�_8H��|��E/%z6zP�w)쮁��R�nzc*�:�݅Ȓ����[Ѫ��?p�Ur)�F t��-�MRp�wh\u�Tw��c�ݾH��9�&��D�`;�B��5Z��
!h�~�=���8E��Gx�E�=ՒN+�'f��.�ӛ�(=����cg%y��	�C��=/����ַ�J����I�s���l�u����&maಜ��aI�(�#`i�1����[� �>-C��ޭ��GP�	r��9��'��z�VtFQjBZ��f�U5ʐ�y��a�#`��,�#�ӌ����sE�'�kL��Tϑ"�9���RRquo��=�#��O�T�<��ż��� �i���ϰ]�UXgR64��[)iWF�Ֆ�A����TX�/cB�:x(�h�I�����R�^ݟ-�T
�q��X�]=��3�V�d5-k����\ʼ��N[�&�����o�<youE��o��J��+�|���7+H��&�'����w+��߾aY9R&�����e�̧������'���u��a�^ ڑ�oT¿nC���`F*�N?��q�H�5H�E���B�"bbL��r�9^)�R.��W��/4�q�s��� �������Fs}[@�>Üo�{*�93�՝�ٟ�F��P7�!�WR���r�g�YnP��O}��5ϑ *vM��L6��.��� ��?־�>�Fy��n���Hԍ�%����E�,�i�愸��+
,w�)����$��Wn�*�@vn��ώ���E�^u7׻���(����ʆ�f<����9��!�u�$�,t?L��H5���@LQw�/_�q{$�,�]���� ,��=�����k��[�;TV� U�&y�����RS�:UI� �M*�N+1H 0
Җ���Ҟ:/kk���Ǡ�%�k랬Fm�y�p�7;^��Q~q�֫q�l��?���� ��e�AW�w�V1Uy�O����n�B�U�Qo���H~�-_�5��:��
�;7�����{6�7=��h���R��*BBK�Up;�w&C�Z��	�T7ñ�����E�|'^걸!)�{=���L��$����p%2x����\��r�����{�䝗�;v�zo��D��=�&��nC(\�dQ����& ��+	A��&��A���Z�]�Q���-3��pԃ����ry������Q��������R�O����+�%Du쏡�?51����U��\샛V;���vq��)��?Y
}��Q+��eZF�l21����b.��4�L���L��ۂyl�b�u`g����ΰB8O]�9����r2pڄ�.]l-��~�ɎnQ��^$���EF�;ay��#/;��Gc�^=#���wj���F���88������BSJ�L�VhŜ�iQ�W>��,V�*��+K=ő���r܊�؎︉J��E$7��-@: 
�
���I)�p��#�>R˥�\��wkO��\;S���DC�ꑙ�T�g?��tuf"~���vv��(GQ��ŕ�&Nr�>������4�/O����������^R\un�4~���70ñ����|�&}�ׯ{`�?� ��JJ�D��f�a#�H�B��5�3 �H�%n�����c�%���J6o]	�x��vy]-��-�S�n�6E�n*=7�
��[��v5{Wg��1^}�����"��,,��2c����oQ��k�tI�����K��l���[�̭��*弓5�b��Q�C�E]Ve����t��e��!�:@�qڲ��HL���B�`�]?��4MJ���d�m���Z<Lj��J�OT�0I���Y�>,�s�����h�k]�q>���
��|\Æ����b��� ����RB�&H����pdsH�[����!��c������`�oE=,�����S�`Ѥ5�#��@L{��2�w��"E�����Ŗn���T�t�}��D�����2Q���N��nb���c�,\�rnXOk�q��3�c  ��+��p[B�^F���" �/�F�����M'�A�e�!�.�3�����~`����Lf�oҼ	�����ń�i7�1R�(�|P�"�X/����4S��ݼΖ�F0A�b����^��6��b��m�Bv��pQ?U��ԫ,�鲠%<)�i���w�eY��e�`5�6�'h�k�٦���3Vt�yi����l[�w�IHA�x� �Ҥ�v;[F��O�������-So�ѫiR�'mI�k���I.�[�;�XV���(��K+w��iv�A�������~���l�q�6x���B�B������2g$�E�ȱ���)̯E�1pQ�I�.�o��fO�o�؀������wmJ�ݑ�hb@�1������٫��S�7�21O�lqx['���z��f��0��^��f(=+^3;c+�Jj;L�el��e��%���A�H��c�U��Xr�Q(�6��T͒�n|٤�Fx���V�^p�����֟`FO���Gh�8� ���֌޲6��\/���t��i)���b�*W���Y�Q�'\NyO��zdfK���m@��Ȕ�&j,�RB,S����I3��J�B#փ������H(�o�y �as�^�-�y��x(۱�b�{##W�gmf-�E,��`^�pl�o�Rܺ����#v�㸿�l�<�Sp�MekjY�bm�2km_V#�+$���K������X�aV��%*��q�ɀ�[^M�ɒ������@�2��d%9����ɴ����K7)��%�"^6}:���K���촑'���
��I�%�`��$Ș�E֋0̅^G�ک���0Կ�힂'6�h�8���e3�-[���'e^���N��	��@�Q�'�*���x����<Ka&Q�e��L�qqK����� }���`�1H���}��	�Go��
��lh�	�OF �ӂ�gS��N}��z	��D�D�T<�}�5,�?ˀ�˹����L2����J�\� �+d��B�,/N�
��� �l������X^D��ZZU���:���oV��to
J�ك�Gy6�?��C<�Ė�e������
{r��n�+lAh��Y��$�Ȉf%5�4�>�9t�Jx8��)��
|�k��.�hbJR�zQ �tq��J�6S��;�!�§xS�<8�8�?#�4=�-��iB(�m-'��E;��Yݘ�EJ[)p���9�u��C�cF�!ߩ}��}Ҝ<V��v�P�M�B�F������]��٨gD�x6$�#k�4)BR�ǣ��8��;����!4�e�tU78�Q/���[OF��XfD�7,�E-���=)�U�^�X�����5���^~F�V�f;2���ٸ�5PC.����!zr`E��;��l([��Ou|�YSE�' �Gy�'��5hr�m���7)�u�1�Tox5���|�z���UU�JT�'����{��r�?<>��>�`�³i}�5��ڤ�V���{�z4�zX Y�.g�U|��qS_�;��8�i\ߜ;}�tG�TA�h�bخo(�W�R�S-��������r���o>r��Wjm�����x��9'����ukE1]�&�f�'~� ɤ�4\��U�#�޻1��e�hQ��gu�ϼp�1ŘQ���JAh�xk[]\��ЌeKc5N���u���rחɖj��]|�S/����a��f:�J��j�w��E�Q-!��v�6�'�*�F��8Cn�.�$�^",S�}Z��ҤٓS�v�
������i�8����	A���IW2���Rn�l��|j՜`��[6o��2B��f'**t�O���`��4�C_�����ͿS�nw$�<�?����?�?�oW��.#b��2��E�M��ћ�5�%W�����H2��{��I���K��ӓ���r�1�l�hۤ����\V����@�뙇9$_������Y�0��\A6D���D�q�J0bq�+�*dEc��D�a5�z���3�.��y2C�?)�H�l�o�&},_钃@&,�Ԥ��>����Mbz�7��R�>˨ZM��UM���U�,�ߖ�Z���͏�0>Op������:��ʞ���ѢO�LV���-1������6�����|�5.�Y@�����2#���]��?L��P�ϊ��l�
���!8�s�M�+r��H�%Q��_=��ymq�ݔ��
1��q.�}�h�ҧ���܎�� ѫr� s��o�x��ݝ����w	��:���,勾���!}���wԌp�����a�����\�����Vh���=�<�ퟥ����!��;QS���Z��(��V�nEA�#�4����� 
���P��`B����m��M�Q���/QY;��C=��!2�T7*El�n6��K�~	P������P� ?�#�պQ�QX��ϱ�A��Ypo&��C������9"9�V�1��-F�kg*ޱ����'���B;=�1����t�g9���l�L��D�9TA��>��E�f�i�{��bw��������`z��G�����w���h�M�<�tNZ�7���m[�a��.����VG���o�D.INٓk�Fʩ!���^�%�~�L��l_�pR�|���d�,��+X�;Њu�H�e	KP_]'��tĪ��4�z4�2�Gq�p�m-��bl�:����t¶�@3��}�ጚ�uA���O��&П0yR-�^�H:�z%!=�V�Cur�'W�ˆ ��M�������bױ�Uu���Vb��
X9V��4:�M���p�8��	�]��N�Dd���g��ѼU����6`�o�v�`[g�X1`@i���ˬǗ�-�>��ɞ��?v�F��M�����4�c?�� �tH.�Or�,�tvc*p�6/< 'x��u��s6W�\���F���?��+��LܨU�{!�R�ED�syT�t�g�[��9�� ᯀ�p�N�g��>���G����v
[\{98=sk%�l3�I���p����,^H�P�2/fCyy���&�w7y�
T?=���PK7�_��q@�f��{��2���0j� '�â�]��w��|�k`WPǔ]_#ԢMzn����J��X��y`)L�<(eg`n����vČi��<:#�0+���b�~�8<����C�_Cڸ�z�)�\����U1�&���^ǺH>$"�l[;���J<óhӼ	Mt��(�(��>{�w=h ��3��r�c,�	=���u�vU�� yK( ���ѱ�W��Gg�.�ٲdǓ�����56���Y�wC��yY3���@�!{�dw� *��QP����z:�t<�eڥ��-o`[�8e�Y:����op���vK��i:���34���r	�b�]����W.ۚ���ٳF� ZW^-��1��̔����7r�DSS�¸$.8K��v�?r��yl'�0������Y��n8+w>{��a]��x�'n�Vo�g�_���H]���7��i2ȻS�=�L�p�AG~��H�N�s����k�fC4u��>��G{R�+bTB�f���Y:+��ݎFtc+��Jjr�����)6�w�����@Ԡ�d=Aln��[U�A�J<=qP�&��i��SW���5̼�s������h6M�$�)|�MtlҀ��f��ޛ<��Ϫ?+7a��Dޙ�ʤm��*)\��#V�%{MV]p�ӱ��<�0=ݛ�)1L����'Nj�q�����%iS��ZM%��)�B��Z.�F�݁��ݔߟ�AUt`��Y[�����Y��>�1�&�t7
|����-K�?�g��|i P*�(�p�6l8�X�����r���<ϵ����Y�s���O��f��#��"_�C�j�s�%I[&��H�Ͳt�:Foj�^3w�����Ol���BK�z����e���a\�8�.�Zl��`CB�#��wZ�)���K�̚F:��٨+Ơ�B?�ף��˫���z��t�0t�b�t����ob��*��x-b�6nc�vt5����������G���y���n��2.S��4�ӳ���ZE�2���}�i�H^�+7�6w�> �¢�l�.�d`/\�}L�X*$cCQ�nK��a�JBjj;L�'R[b��!*�Q�.���(5u=pd������}��_���{�e eHԝ)���#r{�塒�𐐆U"�^���86h�"^���q٦�P$����#ED��c�K������Y���b����C��t�K�Ȉ�Pk'�B�3�"�Ǩ���rR��-�U��o!Ӆ�1R���)�_#�rX9�ƈ��uCb��ƞŴ�nv�x9�L[�j�|c {��-4�݃�������?4Ǚks�k�������D#@dę@5��g���q��c�hw�F���R��ݨ�H���m�7��r3����zw��	�'2e�o�V���k���+�����S֎Qt�t�¹5���pc\/���"ί�б39w���c�h��)A[����������� �Iw��Vv%8����Č���Ӭ�M̣zig �(2�� v�������+��s6�g�Є�O|��k�Ds�{�,�2�V��s�waۯ����K^?z=��,둏�{�A��Y<36#yX���*���P����d
�w�ĹN����%hͱ�n�)z�(��J	�����Ui������\��ڳ2���	}0�焔��6�(��j�h#��OT��	�7;�3o�r�`��7��O����Dݤ���q�ڄ��-�'�L�b�UsQz@:A���,�aV�.��w=�to���.�l,�iF�����حa��tG]�`ru�6F%o5pn���#�ub��I9arD2���T��W�C��e�]�����}���n0�&VCp�z�$k��G�W�$�.2<�?Z�(d�Z[g�"t���.:��c�f�z��K�3|�yٸ�{�ėF�	zi[|� 熯��P�R9��Ej�����sn
k�X�.ڶ����HC�	�K�L�ǽ&��'���=5BM�@�3[^�8��-q����q��D?�k����~LmC��Fl��\L{�lI�;l�@���V�Z��,?'�QeA/��ְ����k������������7� 踨����n4�<�2��sS ͦ�}�����\�����Z�I&�Y�Q" ��N޺���_g��,'��vA�����W�x�מuYr���,u���Si��B�1�JG^�e�-,M9X9���������8�Ъw6� g�c	(��7����2.�An���3\T�U��I���z0c�[g��q�NI-�ѡ���1�a�c��Y��d�.�� �!0	P�F}Fj%G���́i�����r��,��[M����ߎJh9��^�V�(Uq��	`�8L
l|"�q�/B5]1!�7*�:q$�Akr'!zY=��� 
1���u���K$�
�ǫo�ꊠ&U:QG�����k�j�˩���yIe��z
�f)����A_��G8X����EtjcqQZ��f��4:h�{�X�t}����kHF�[�g���4����vW�#H���D7F�zx�S�'[ ����G�\Mt����nEV������h0=��<���Xk�b4��t���-�* >X�Sl4�	���&8���b�"S2�G�,գI`�h�}T)[�z��
�6\Y�$@!Έ���V�l���cKH���ph�7#�.۫~i��WE��T`z����R�U������T�1)jY$[�U����7�#Ӏ����=��kn�)�@m���ܩ7t� ���X$g�ke#IN����Jx�BƠ�0��B�օu%z$e-��ؐAQ!*�;L#tS��!��r\� A^uo�E/}e����ie0~�q���ѯ7���7A���#+9�Cb�>i����#�K%,��"��kV�O$/��{�RMγ����Î����+���?*��n�p�Km�Ly�(,�:��-��q �
�H
�PZ9��讱����`��ә:Py�)�o;��~��	)�R�L����2[�#��J��۹_1�fO��_��8孾/4�%�w��������?h EOQ;	�q�i��phdf�Ojl��bv�i������`ci��h�:Au�6�R�DUBC���B	l[�9�˰��(����)����y�EI���	���n`�$�	C������V�p]� �3��8�RY�,��e�6�A�/���E��n�����m�۴�d���<�_�J��	�[g���N �#I�͊nZ�X�pM�t[\� 6��6�<��H�~�CG�$h��ss��0�X�Dn��B)]ԟ�f��Hkw��O�^�I�\�t����h+�68D&��z�,�G_�j]�@M�(n-W�Z�8�X�T��%aD��,��tW���<.�8�إ.����8���lzˮ�ۓ��U�	���ڎ0���6
�K#~<���iGLRu2Qz��N�l����A�U�X:_��3ƌ{���m���!G����]}d�A�o2o8�_zy�+{��Д$�����%/T�C�gH�FT����q*����FG��v���<���"���w=����&@�tϟ�!0��F9��M����cq�?%)t�|��\
�?��o#��t�
�	�	�Jn#ui�%F /V�������-ؿ̤hk����.��ʺ@A��+<;�u&�8�$��)��6|�����V�ſd_Y����q����(w~��e��j�zL��t������QP���j�U�P�"_a�e��G��`����GC�vt&�4�+��2u�"��qpC-P���.��M��, o�2�ײ�����.Oݳ��e�W�F����_�������:t�5���{>t�����+e��$>���I�UNz�o����e{|;��8��[�0����;k�D�p�g�6��a���4ߙ�t�G�2{&������lZ�c�̡�&|�͉A��i���5�b���%�zV����H�[�Ϊ�&�D�Z�r5���x�]
΂=y�[F�������ߴE�ER�^��@m����'w^��o+��1���x�^xY�f%
7S/�����?]G:��}��=�X�q�R�cU:�ݛm0_��ӱ�N�ѿ�^�H���mj��� l_�7?��"�V3���מ�8��޻�8P7x!����é�?�G�҈z9�Ņǉ����a&��h�ڸ~���lz��_gyu<���fxx&�碊���m��rZ���J���Q�E�+:�H�Y��ͼa����}Ζ&§����������KO�x&�T�޼~eo0�d��bPq;�>~�G��?�3���N��1��*l�'����q�*T���u��d�/��kC�X�Eo鷱F��`��,�A��fh	C��S4�/�Qؿ���A��d��5y�A5�1o}���Mv��`�ׇ��#�Ї��'QISlp�-��U��ҷ>檲��ê<_.��QPnV9��1�{dK��
^0찌��ش`Z(���1lM�v�$��7R7�<���r� )�)\�{#@$t�8[�*D<�L���� Ԕ*	�h۸��G�;a /Ç�mg�>��@�wtp��j��Ѻ��Y��"��J"��2�+y.J������U]��!ta���~��S�v�M�4����ŭ���G���Z�&Zc|�y��O(c2?��okbS�.$�J8�77C���qVA�O�p2�꧓�SC��wP��Le\�� ���$�K��$�4����Cz��O��-������a`�Ϲ���6o�ڙ�b.��4����\�]u������c9�
Z��C��{hjAPH�\|�k�h�F����!1a�(N��0al:����B}� G����Ȓ���S�s&�6%W֍GJ-'Z:ɹ*�\ā�tX����ɢj������Ҧ�PJYdLxx�`��>�6y�ڼ��a�z�[�������v4X|Z�J��\�5,�I\��r�>���pw����76�S�Y�eZ�a9:�����zA1
U��Ĵ�%O���4��,�Dш;� %�]���@Z�5�4��d�B�hMy'�����~�I�THS�P�bI��:X�eK[\�l��+wb`��p��T���t�h��O���?HA6�Q�*]:O��¤�}������������\��]�K"� �l��$� �
O}��`ƌ���H�z�n�9���Gl��>]i�)ði�(=&�>�C�	y�B�m�����y1���*3J`����]�5��J[ƹ�8���� �}�
��;�ip�gg2�Ix�r`k�da�o;a_���[����J�K�g#+ךB�(���j �	f1_�b{���!��,�_�@��FfEO蹔*�Ӱ�o	�҄͹�|�K���ڄ�o��dȄM ��kH%�J8%�ٙ�4��	��j��b�C���4F�S�RY,��:މ����ń�<��^,�o�Hጻ�xD�\|¦�M���Pi|����3������j�3- 0bs�.*�(������PghM�|��\�T|�𱷪j����6c�N��YS�a畫=�m>4�P�����_?��wf&�IP"Y4���6q S�L�4j�!���qH)&��j4'.�H�VU�������V���q�� &\/a�{t����3>����)ړ;h�d�����"b�soC�=���6<mk�%�\l�q)"�.g����p#��IĿ�Fy�f#*K�?�>Х�(���Ni����P��l�P/��hN(�#OJ�V�ݚ��	�t1	���q&��*��DN�>:�y��ގ)��?(��"�O,��A]T�P���+d���9������(JⓅX���)Y�;?��� ��[�F�� �RCe�&�Ib[lk\�Q��;�V��"��)�n�>)�G�~7S@ r�4Q1wJ�!�T� ��@w>��#�61�2pQ�O������� �ܬ��Lda"�د�>��c����=�!*�}�W��$�c[WYB�M�]f-_�HCZ=˯����ѱ�K�Y����4<��Ԫ��^d�iי>������k�}6�2�1p8��w��#�+��� �,YsV)�,���@8�݅��}<[���k]t�=���n����*5�I	!
���|$OL1��l+��V�-q\J����FpH��f���S���4�B�xI�3"D��FS-�W?�)u���@�g���7  no��)a��c�A��MSz�Z���~!ހ28�>'z����qX4���)�,����~��&Stb�-P�����=�$٢���g�ܑ�b/�E�\PFD!#Uf�r^�ɬ�a:HO�x�|R��):g�	E�'Q�DX�]]�<Aŗ�5��B��ź��]@>�"���WC�h����0�,��}q�۝@E5`��)1�:�//��6tA�qCސ;��	Íg������T�Q�u���(L�c��
��Q����Q}�I�)@c�:��;��x�cUܾӿ��x�+�H��� 	��뚥'�|
��5���ٴ-�j8��1X����K�9�n�ܵ͌�H���Ū�&(B�d+B���u8�QQ���Md�"1ڻ7ڷDy�\Q�����WL2:٬�m�,��/������I}n�=���6�{�'�����n��RH"v����f�^�����:��E2�L��t.�"�_��ҕ��/څݰ�[V��5wS(�Z��MdL!)Q�3������?j��犁P�-Mz X,a�3�&-�i�m����QR`8YE3��h���%���YM���0I���l�+��1�E����_��摊�}q�BǤ�i���u?�E����ȁ���ܑ��ny���RFo����� �=?�R!�٤J9(kJ6���	�������NG�t6/Z���k?brC�8�B�˱ɵ��x�0;8�>� {5K�x�eǪ;�V���~�xBT���Ʌ�|>Ԏw<�n�)�4s�^�҄ VKq�1���D���݅��d)%�^��ȟ1�đ���Ku��K���cG#u��ڐy�����;��/a���4���V��x�/��#cX�1�׈���� �f.x����WA���k�W��c��*r	��ٓ�XX���:nM��\9��`���(�A�̣2�)�G%&�H�DO����>o�iȠ�<��MnܞD7W_0Kĭ��8g��$�n����(��`�T�n�cb�El!d{{���p�W�w���@���?�S,����\���������7o�����7,g��`��ʕu}U�.;�k=�=���QR����W����	Y�e�ɶ��F�s�H.;]��)1����I`w�E���ӏ����+>l@�B��SܞDad��	qM�>7zl/��Ey}��?͏���Gu�0<�ex��Z.[�f����@!h�u	x}������O�s,/��v���U~Hg��2x��>$��4��.ʠ���BgP��z�dQ&£K((�rRA>���>n�l�H\�������}�xIP'?wΎ[�Ǝ�n�6���6c��W��G�(�,�o���-��n"�mܥl�n�,���ݔpޟ7����#�"��-a�@0���`pS��=;j��>u�A^VaV�����&�c<B����{��N�ΨRa�X	Z�g��R���4�Ι���%�E8�Q�� �C^���DkE܁5�"v`�ݾH_~�.��4��8>+�ѓ~{�%�m����,�c	��{s�����74q?�G�E�?���[l��t	���b��^jc�zo9,lj��@���챎R�b�\�ʁ��`�)OUF �q����=~$�q�P�2��CtC��/eʋq�����>��y�~W32^��<4(ݍ��8s��N���0�L�}f^��x@m_��O����G�s���*��ǮQG/3T��2qoѣܖ�ަD�mڦSG���ȈM��Z������t�>��﶐�R릵S�����a�x$Gb�><�����f�<N��qX�m:��-�[�W�Ĵ�t���=Շ�Iy#���0���5AkXk�@@�$n���mh9���z�z{�d�ٗQA�{�ʾ�GB������αVu
�*v�����鞧�9��b���%�|����ĺ�;��ּ�Q��"��B5� ��N��	zO��0�iW� {V����)葪\GXk]�0F�.T/ЕzV�/��*��U�M^��;��B���3���)�e��H��_��R$f�[�}>����8��eh�A���4 Q*�1֧����!���h���(�o�N�0bW]%�mfH_�I���0������Mw��+��A@gl�"t�W�7kذd��<�#��=�U����}��V��VG}u���!Tc�׃T���3�NiL��sS�ͭ�UY 3ѐ��� �����{߾&h�%ϟ������l�8:
�o*�0'���O�*A�1��_�]g�i�ƭ�VH=�r���e6z�#�b����rZ��HW�R�WP+6�9�h���>W�O�n�+�g��������K��������~da��y���XGO�?�Y��e�ݸ��p���H0v�K���7&ʿ�/��:����*�ǫ8հ�Q_���|e���?2��Ix��Ԑ�Y�2P�Mw�R-Ԕj��b�eZ��敏�a�$w@(E*�:��i	X�5��(^�@�3�+��rz��zLR���WWE4[��U�	I�2p�t��k8�z�0�W��K(YL����vS��~>��I�S���v_C������%pp*�BMm	k�Z�-�e��y�Y�j[�D�U���_Z�5����.�"�V�?�+�šr�$#�!�K}3����<�W�l�4�})pQDm?���K�S>��l��Ii ��ސ>1�,��@kH̿gP#V���DK�u	�5�2>�`!&�Ӄ/��+�_k���'�	�7
�eg�E�d�m�������w��x��.��]�r�rH��Otƪ�gɼKl�~�-�"��k�XU_k�������/,�B�n~j�n)�y�Z?.�/o	���A �Z�]I�Mx#0y��r��5M���'�����E	�-	q_���"��Sjih!@���g"�U��<���F3�K��Ch�d�"��U��å*�����:�ojN��xy{�Q�����館XY����*n;�(��!�R�5�w��,���)�Q��3C���<�ų�^�Δ��7J#7Y�ԫp)桞G���_��,��31��eU��`f���k^� c�6l�x�q�qZD�N�C0[j��mG���Y���嗽f���4�����h��dj/8�E�D�=���΍�V9>:Yv�9����u��N�-���:>����M<x:4�̳$���yn�ϸH	w��C��STi�I�;�[3W�u�cm��P����|jUP�w�o��˱q���GyB.pequC�hг�C{��)7h��xX�7Q�3�!��+�/w&02r?=�wp\s-��I�yc�j���W2-W��{�6�=PL=TY������|�.��h�=�a�~]�<���z���cd$�xd?Ţǔ����wY/����|����������4.ea�I7f�PNƠi��A�|����"���𘗞JB}�����lb-��Ѱ�֕ +b����V�8��v�]܎�z� �"l�"�%�Rm�N�vLZK�!��ܚ\@R�{��7[�z
W�XS� �A)Jx?��V��~μ��/OFt%��L���3��e���U��F�쏐E`���x��ԏ����ӀxS�`�m���jm�h�J��NZq�h_���J^��x�k7�p�L���]`}g�)�׭�ӜK v����l�d���7��6����J,�@�ͤ`M��/�QU|_Cz�c���������#����4}%�t�o s2���ݿ�������j,�n�mj��|��07��Z请�Ƭ��Wg��}]�J�_K��򆅋GK�	��v�	������|��3�C����Gv���%�S\�;�#�23�P�_�3:���@�}����4>����c����ނI�g|IT)���*;
�PQ�a�/�aۙ�ci�����	�ծ4!0ұ��a����H�TLY'��S;\��ǥ��!��+bշp힌Nh���֤���O�J�SQm�I�~$�Ԁ����L�o�9X~OI�	γb�S�%�ɛ���OD�ҷ<@�ε�\`�Ss4ŰY>E��f1Q��=F�%�{g{�5�8�y�/�0�;�/O�QC�8�D�E*�;	Ƽ�lk�Nǒ�(�����7��s[)7佮dm�$(Jn�=��\OۑT�=�a������Ŵn�^�;�J��T��5�����	$��{`.�y�ν�br���5���f�� ����=�9>�� ��R��'���<��#KD�9f���DG��|-F�wL����溇`�F��2 ��5�h�����|��)g�� �?|�ف�6��J= a\Hr�Rx��!�%,����>7��}��T��5�'XE|EFw�G��[����c���酶<q��@�Z
TS�1�ɯ����u�d[�_zW��̈́��7F���?��1h�8AK��ƺ������R9V>	(������Ԇ��H�m� ���C_A��"O�c���l�cyio
��ՓC�vn�u'n%���0*�����E���uv�6��Ňc}U���%G4��tG4ō/h1�Fn^9�W����yb_�3aف���C"�y"{GO��(=li8���{����|Gml8������9w���B'wM���RM��w3�܉s�2`��S���,�'Yc�;��%�G����B�`�a:l���Ͽ�o	������q�o����2d�W������q�d���wz��������
�9�Tj��J���R���&;-t����������ےW�kXi���y3x��(�	S�uT�Ǳ�}�Vo�*�i�����&���8��m|�Km�n�$U_�?�9"��)X������i�o�[�(��и�G==�j�P�/�Bf��m�Z�2�ړ�L8��f�I}���x0�m3�fc&��R��"���X
0�������ΛRth�wm#�8-�m��C��̋� ��*X��/=!쫲Mr��In
�q�&�����Z�k%l�\���A����|�=ֶ�|e(�4MN ʦ��q�2ߺ"K��6�������T��>���u���Y�Kz��Š�!+��1���9�[��~PD�r�z��$�,�G��?�x!`�Rʤ��fe�<�p�p�����&;X!�����y����۷�@���$o*��G4&�q��k�TZ���/���	���ͽ���@�_����[�� 験�to�Ɏ��f�}=��w���3��y]�sN/��L�	�����1��B4wm�6�l<f��"n�=�?so��#�sqQctnQ�#�3�ə�$e����D�T.��E"��H��gmM���}wۃK{ɑ��Z"�,���J���1U�᝝������]�u�CI$Rm\��ǟ���,�P�>9�{�]'����Q\L2�����$��K��ZڢP�2c�@iǟ�;S?���z1���t��vU�e��;g��%���':ِ>�\��fP����}BNS��J���s�y��ÅصJ�Jӓѷ�u�6{5�.�R��Q�W���V|&#۽H�X�ʖ�!�[E8g� ����譓dm፺i�����8�"�r��/��W^��Z��7��B>��4ӶM#�t�l᷆Q�8�{o���2W�)��ߎ��		E+�����n�Փ� ]�r�%N�0��U�]&/��$û)j��e�ӧ���@�,���!�\���)~VЧ�՜vƢ��+��A�� �@}J�����4D�O�֕��������*ؾ�Oho�=%�<����Ǉ�D��_��������{�3(��'k�b����1*:A6���/���M�I�#�8͹� )�t�uirO|1�p1��Rk�_M՚��j_��$=��E����X�Y�0��EZ�:�~���g�qf*ۥ��A��w�?E^���7�����JM 7����u�&Y���%��n��z�S�qY6�k��,��)��hX��O>ڶ��F?����T~|��F�6�y����8AZl���ZO�Zx��`Dȷ�l�o2��9���ǐ��>ꦞy@�؅y��f2�q���w����C\Ĝmvh`8�G�[B�p��T;�����r��y��䒦7��v�e��3Т^�8��BZ�C�m�L6
��_)@-�*}�ݔ����ȴ} PF��]�����	�ov�&��s�<0w6����"����������Kam�O�;$�ֻ��(H�R���m��NT˭�܆l��m�d���r��yv�#��.ڞ�5Lzli�%�P�.Ti�P��[�����5�ǋ��T?`;��l�Nfv�7M���|
��� ��O+��l�� ��	�!�M�/�0u�RWu䶳fr\�=fS���9�T�c�6b�X,�u٨v�����L�	�4�P�Pʝ{_��s,��b�إ��[ۓ$�T��O���j�a�n���?2	���%�@;��$0�n	� g@�����gJq%�N������RP6RR	J����Jstͩ�43;$�cm�:9-����4Pd��B�	�V1���}��	�å�gJ ��^���Ü��ϸH_2������y������#�����X��K��\�^F�e�{��e �_�A��i��%h�u4U�Oy�l���d����ۥ7є�_�G�ߞ�E�$V����������^:�)��"_����:ᡯ9��N�/�Zn�cnNf�r��n\��I�E>����]s
�rk����X���D�?��0�y1��DNة$/�2NgR�$���F/� ��`KB�w$v��^�枟�/��6+�4|M�Ʈ�O��ݏ���1�7| It�� �Ywp�%�i
��j��a�Hf�0��tiv�粅�/��B=���b�#H�Q��~�g��Q!�%��V�z���t�[={~K���x�1�����+4���=`GJa��n�{�7>��yF��8��j��g�t��@�5�B}�e���g�\��y��,t��1�
	���8e_�7�_|�ᎇ[ʊ�q7�N�'�֙F=ɒ<N��8�-�V��Ok
0f(k�hf�t�z�@=#OJ���������`I�E;xf��:�����Ϧ~�����c���ӁDah�xݸ�Cg�"4?4M�8˨q��[�#��2ޠZ������8�h~ܰ� ����
�D�{���鵻�)�b�6�d/e"5뗤/�d1�)|�ǴW8�#�w����g�x��k� �6�Bq�EUc0�`��}K��i��<��^|�4�O��1^s���2؟M�>�鏆.�K��\�'�>����Q�Մ��b����Im��"���5��SVL��7��7x�ȳ�X�&ܯ�f��E����f��Ъ��h�vOS�����}��|�ם��+�~�Z[�.?D�(��h!"a�d1W_1DBE��<2٭�Fb@��=��ԓ-[���n�T��n�3`%KFB�G
>s>�R�� ��YpEM��i�����=��/��h������Q�?�5'�B�p���IY�}�����V�!��=cVn�f-]��	YT��#�̀ф��5p�����B�f��ۂN�5_A)����KQ�0�ud��m4k��9�E���l�iG�p���t�����a��u���o�p$�4�Nɺ����a��T�-� ��>4��k��~�B�BaF?�� �����#��i������ޜ�dg����8$=l��R�|�lM�vc���ZЧ����[�$�'[�(@N�K����!d�cb8�M(��f;�cn
���������h1��o���ö��H���)�$/-�18��I؆̂� H��G�S/`I��@H��$���?؏���֨�ʐbJ)�;�l9}�W}wN@ys�`���&�Nޕ�)�S��QD�ǈ��!��0��ao���ki0�Q��ƍl��z-hA�Ӷn?CՀ��U��{�CN��P�<��r[��5vՌƖ�B*��*����zsl��� pm���h�g��I�% 7��Jz�5z{#?zd���Y�UR��S��a��]>|��_�5��Pځ�������.XT-����5݂<�7A���ONF�;$�b6�&=Ї�V���R�i�[�����~}���PTC\h4%B��Y�O����kN��FM���J���\T;���*̰�N�����(���7(��llC��4,��^�Йʍ�Aƥ�#��;���r�H��P��aR��[��F�=�E?S��?��MY*�ER阼y'������u���*׌����A
���0�J�\5�g��{-�n��R�x��A�P �|��_�����"��i�s�Nz�W딙v���0�6��q*I���}t7w�[T��|��d�V]�J��n�kh�Z�
BD5��,�)M��G�7�y��W�y��֯��9�¼Y��ä�d_���S�~͊l%�O"�S	\0�bC��:)B��2"��9��ۖ���Y�F}@l���7ifn��8Ѐ.�|}PI�����:�۞Ƞ�2F�"/�j#�>VZ+ZTCI�mx��o��x��B�xұ$;:�A�)^Y�jL�����v�g��Nݻ���s�#�:�C�%Iy�ll��~o6yC=��������{y@�:�Y�J�AP�u�zi1~)s0^����)��9Ck{�(#�K��S7��#�R��=��z��a�=1�(o�r�{�!ή�hd��+Ds�=%{��&}w]iV>|�x����x
�L����+/P�;���ax.�P�9����\�b�J��A�{:�F��+Hj�8��	�AC^v���Y.A��\���z�{b�����Ř
�������"�?RF�V5��x�����xZ��}ߩI�+���E��D��vd2\�^7`�2��GeNE��+����p�!J-��4Zk3�`9�'�j�P>�^��)�$�:,V�� ��h�f:?�\)xh��oʿ�ǩ�����%�\%j�U���/3`T�Ze�]R.Z}J!�Wc+W��{<3p��"���X�qs�!���c�?��!6����{V\oY�Zˣ�{����zd%fGž&{W���{<�ݡh>k�6�cܧ�(�:�����n��O�L+���t�Y�m��}�?쎫�9bs�-�:���Txs�̪,�(ے��p�[�;'�G�Nv ��{��zP�ܺ s�k6��6=�)��Zb��=f�~�J'�L��6K �*�� YIa)oK��UF��ӑa��
�!��3%�RP�ͧ;}*�+S8R�H6�i��_����`.�9RN�V)»)\Ǘn��]9� a�c�Z���?G��ȅ^h<|�սΉ�ߏ��3V�Y](� ԧ��է'peW�������+Q�!e�^r�':.w�,(�ޭ��S�Q.I	�%x}:rE��%N��U|����Sɻ���誃��"��$��>g�[�MKY�V*�5G�g�%�j��k*4-��(B���o�������7P�e�7�]ZW�hdPd��������*��T���ׇ����3�(�eq����N�l�c��}�Б܆"�B}���c���xdXtd	)�R���}���gVD\��o�E�LD,�ױD_���Y��b�3_�sJ����b����ڱY?���X��`D��<�̫S��E���^)�ve�K�{dG�+��gzp�NlQl(L���4����$�nB`S�/X���V�^u�i�qo#q ��D$	�7p*ҷeV��5< �/�^+�4(8�!�x�H!��u(FN�[���ގO�C/;{�5�` �]�:����EP,Hq�x����;]BАA{`9%	1����F0:>��5aiK7������`��7F��L��3�?:~s��@4�M��՘=}�?�N�������b���UE�����������m%���p���s���,-ʆQ��⛆&pB��%���в����IN]��ڰ������Y�_��IWR��+�-F��-���������l\�n{]�8�!��{�V���2�z]iYA}�"#�u�SJ���74��d��<���r.Տ^�).a�g�RFr���e-$�$(Y���G�Χc�xR�v4����� Wᑾ�&��j@=P����h�;���88w  ~�J��0!�gd!�^2�E�;qf�2���m�W@YW���i���$^��K�d}��a0��嬆���h�Z�"��q�PՏ�)*�pʕ!�Nu�pld�M0Crs��mP"N�3���:\�~���(�d�S:�{��?�~?���Kv�E�|����:d�ď��*�@�T��b1�-҃�[���Ql�I= ]�����-rƒ&��'g�fc(k�����K�`�jd�/�ӀT��4�����s��Ś�J�0\Kmv�\��68z�T�9oOt^�����H���|���i�]'��	�^}��pC��������W����B���^��z���Z� �q.W��u��)���b�D������=\��l'���`��Q����B"���d�w?_��L	���Ov�����ͳ^s��4lP%E���P��ᇦ2Q�;(��ŷ.�S�� #Q���-�u�����M�1���	2�Z�0WrA�t��I`�u�k���1����$�E��9E
+�?
ǯa��@&�m:�li�޸Ǹ�c�q�SGp>��J-�ޣ�����^ȧ��l��2�,=ʧ�Suj��hP�YӜ_�(Z��>F�/�C�����n����ZN�:�KtDq�N'�`o>]�r�<�{���{�fд9W�I����܆��Q����&�X�.L�<��*���zq?#ˤw�Ȭ��뷌�Hv>�
���Zr�E!��uƴ�\�6k�t������'�F� �S3���a�Ox�����|X[!�~d�������)�)@@�Z�>��©JO~�;�2xN�\L[k���VL�M���6�y6�����m��kY���+-'�D��f1U%�( _��*I�6���@���W���>���P�����;��~���>	d�z2D��5m@��W�ƽ�,\�����h���X�d�_���N궓{���M2���͡��Җ6n��̬�n=	Y���ac�#������*7r�"��g��f&-d�2Xă�497���վ �q���Uc��/F ������-���o�gg��V�"ݙ3w��Ce�Y$[�8k� D��$s��|��o��v��RH���m���������xe�Z�͚���*�uL-��9B��צ:+��L߼l�n,V����yK@ ��hBY�Q���>�dh[.[[��dA�����zv�V�5Ӏ�� �C�Z�H�	�%��f4U]�)� �$^��#eڞ]4x�ç�6I^��Sp�NQn־������kV�{;2�C�+H[ce�{o̵f���������I�r���"?w��6�"�Hc����;QSԺ�_z6�3��\�t9-o�&�'��s~)�	�{�n��s��cZ������$�n���lh";��XЭ� �3z���,ǈ)�,.������ڍ��G?BxT`�@^��ං��_���8���90���͹�4�f����jST\�q�^HY���v�0v��U�i���vJ�M�h�]bmvf�'���{� �J~2@���tLf������ �S����9k�=�Ḱ�+��#3u�@i��^E�f�c�Ρ>�q�4ȔЈ����8����]����K�)E�>V�V����Cƙ����:߶���Z��qa��<��6 ��9u�d�[�M�d�*ܔ�Ȫd���?���A$��]:zyy�t�)�Mo�@�����vw��h"�h��:X����f�%����Q.f�����������G��^���Bw�*Eq}I��q� �N	a���p�8�&Н}8Ҋwf�k����<҅�\,�� �y^�<�;�*"j=�p*�m(f�ޱ\�Ɂ����6�9o��z���ř������0��)[�9א�����;*z>��ݧ9�v����o�ZV</�<#Xu�)��G�jN=�:˱��Z�lG���KrҜ/���QcE�I�����
�b�Ƈ�8H��Ll9IyX2�MZ>���o�}�ҠD{����J���bBs響vF�$J��{!ȳ� �x�,��8�����NY��E�cdS�8�u��ǪnRi�{3	�lY����W��0��)���y3_���Ϗ�\{�x�X5�Wq��n*'
����C��C�7���n���C`�9�U��(pj�C�a�Ƞ�bҎ�5���hN�'���c���~�e8E����c�Ie�؟FΈ�
nK�&�w��ݶ�m���/�=�/�M��*r�T�[	/�#�_0�����\�����6~`���ZByN,�z�]^1a��h��n+�6'F��lH�ׇ�x�ހ�+��3�)=��,����U�c����QKV5ꥍ��J��}R��>�ԘE.���Ј��P>�а�j�0��h�U�垿��K�k�Q�s�0e�f�T�����=�EخWP��J�˦�ʂmV�\����(`���g^ ��� w��Ü�����Rw0�k�����_F�M��+X�� �Gs�����ܻ#Y�c����Pk�9�wNsy��(�ԏ�
�����D�5i�UA4 '����3�I������얳�nc��ca��� �ٷS�� �{�+�w�<�EY!��?Oas��W�(G,�"ƥ�����R b�����u�{Q��a��g�ɖ�������F%�L���0g@(ķ�SSA6n�S�?:n0='���0�ih�- Q�au^�n*V��
����L�h%X<�Mi�A�=Za�0!�S�E5k� RH�y)���:�l�N����h��	$ꕎ��ۻ]�<T���ǼzL4�n��y��z��?�\�b�s��F�\ƚ���_)z*�8^��`��ɺ�@�wDc��%�EI��^y��}�O�e����dtC�N�c�S�Фb�iܳ=���z���_�e��޴Te��ۓ�8����ƕ$������`&1��'��oAK�S(��c �-@ٜp�8�J�
u�Fy�}v�ǡ!��M�JfQ��}�2$�M��e�S�C,�/�+�ێ���j��r��d�Լ]*������U-�srW	�����L��j�ED�z���4�s�O���~ �^��8��M
�pѕ�/�?ى⒪�p���kV�+<1FP9��K�����V\"e���[�����ց�v)3J�x�/�WZ�@Qٸ"���|v�pXJ�a)2�c	 �B!\w�GU"[k���X�,ZR$��FJ=���kw���ZȮ�gK�|��&�U^f��xr?�.�uK��'�J���O��0q�v�*�av��c��AR��e@h�B��gԱ��l)���Q!gX|�C2��D��@� Z��2
��H֪i�U�6
ɰ��b�{yR�u��Ԩ��9��6��/"�[	��w��n(Q�
��܊p�$Q��<p�v���#�7�q�Nw�A9�]���ʆ[G�`�(.��m�5�P �w�=���G��]��8}�r��������^!Z�8 ��Q�h���Mfd�"�o�۾m+q���H�a-J(7��}<��6*�8�Uq��P	��G���#�d!�D��K��l�.�e�_�1}�ѱQ���؛���so��9;*<��n��h)X��[`!N;���I!,l2��{D+8�I�S��;��rH7���춴���s9��c�R�,��!��E^�|t�%��UB0)b ZԻˏTv�3����4��Ú�^�a�9���#�ShŰ]i2�WT�GZ�f�$�[5�Pb!���d�dwT/��b �j��ݵt:	��������A7��~&C2�{'H]�����B.i�e�����*�}��Dj�miX�s�'�탔uE�ù�d�"M���nA�r2��BwҴR�e�?{�,�1�Nz���as[�Nl/���[�׊���
�Xg{�$����e·8����`NF%J��K�K��bd�N���T =e	:�<���F�b�����ݧ�'����".#4�Α�e�➣�ـW��N�N@�`լM)ɱ�lWTk
L��>��_���	��	���@g]�?[l]�ǍM��D���\��H]
��R�˺V�6[~�rcM�����y�����������?	��!-��i���f!��-J�����9E]Y�,	Sb`����V��&x�;��axd���\���2cV��S�᲎^/6bz��)�y8$��.�Y?o�
��8�9��fr$.���#��9�Y:YZG�(�����cB��m¸�+����2.^��fmz�)�K�3Y�NGU`H(�Ν�>�m����8P�qTO�s/��𔥲M�Zܥl)��b+`�3������ח�N�t�	4�J�%��|.X����t�����gc��F���~eNgR�	μ_��`q���ߓW5t��)�}��k%ƫҭ��4ȉ朷��/�Jy�]�v��1͛�e��@5�5HT���"31�q�q���:���)�Z���-dku�i��E��vC�Ĵ�ݳ+9�gk��&u�? �C4�=YK�VG�"�LG��ړ�u�]�T�{������];�9y����^
sB�k�5W1R�Xt����/���\j���wi��a�	�+����hg�`9��'{��Y�~�:�
Fd�$m�Ϣ�:�+$�ȋ����-�Z��XD��1���?�+0�Ѐ��GVp�����9[��z�c�%��螭��	����m��a=����gxX�3�>�$��N�GN�k?,�k{MK��Zn ��H�]�S� H�ڞ�|�q��0#v}D��׊J�&��u�&�aS��0*u�$f�����U�p��옿����h��h��T��41�T���Mi��,E��f�鍊2x-
��q������^�9���L#�>�ҿ��4�9��?2�
�B%B�vD����.�Y~�h�4�-朚/ʏZI�	l�����G�E�8��:}4Ф�����#�|܀���R�ؒGZ���~P�ӳ�+����A�bG���[�{��,�$b��#�2r� 4.��c������X�
�q��cH'˓���}�F�D�m��(���(EB���\�1z�7���n��5U=4ҵ�L�oV�'\$�X>�j��+$FA�qJ,YDd��Z���ee�:�Ϙ�����S=�VRS�Օs �3H��c��t*�w��c�*�q�%�����}��=�ti�Ç����\.����,gs�ǟ��YCt%V��d��#�Eb*&��dԱ���t�F	(:�t�Z��p��_{n�J�8G5D-�W<dڡh������oݪOe#�P���M���`%�x��R�H�ϒ��Ԃ�6yh; o���*��ܯ8�A�n��s�\�a�ҵ��mC�=,h���� �`-(��}�3mZߊw�L�����@\��v� ��*v�H����kd�xԵ���I=?�z�w�|K�H���Y_�W�� ᪆4cm ���"P�%H��9�|y�߬x�u��M�Ź�#�p\�G �<??y�Tq��f��/��GA?�*/�bL�K,#W���xe�Pksg{����h�
�
�"�胺�n�m��P��o%�X�@�Ɂ�V������s,)*F��5�C��`�yT�����~�NF�MI����r8꺋�䶩|��l�z��-�<� �b�����p<Q�i��&�uw+�}���^�}��k�f���f����ǩ�IW�=ܘ	u�M?cզ#����}G���Z�M=L2D>�U�P������V+��p���.s��������0����tE�YR����{\���(w��Zr��D"����B�W��Ĳ�fס�	��q�L���W�fݲ���ȱ���E�\[[�|�B4�R[�@Cz"�z��p]����k������9�7$]-HEZB���~�ŘH�j����ic&�����*h�z�F><�W��c����$rauih;��9w��<o�n�I�=o�=�+ǮV�B$���N�I��E��ԗ��D������p��C�k�.��a�^���N�A����_�rG��'<�3+���.ڶ�g�u�����2f��
,N�5�Z��F�5u^�v�X�ǪТ�z#��'ke�g!�)oЕ^�EWA������w��!ً���Z).��Ӧ�Ǿ�#���m뷊���ÊK�<�ABz-�:����K����oX{<���tI� &�1�>Ȟ�_&��5�}ˈ����X�)D���.�%�7�.�M���y*[v�	6޿Ů��w�A�4ь���n<S*�����b���������I�D�h,�%lI����s���y�e �:=s��c���*f�Vj���$�<sl�|f�X"�Pg܆��ZL��k`W�����F��3���[\�B ��k�V���K�+�C&��+4;:v%wR\�<��Ҏ��R�ef�_�Â�B50���?�ȻUb��s˺ec2��+F��XS{=w��!ـ:-_�N��>i.L:��o�j+��^�5�#x�7s�@�IM��ܧk
b��^�܄���*�����o�3�����Td8#��i�<M-K_�Q�&4�w<�V8��6�v��g!��޹�=�SjGF�.��vc�ɴХ�c�/��֞��(E�����_?4ۖ_�ԋ2� ��`%zC�s�Z�g��;*[��sk��Y s�aU�4�o�D%Wz*������nZ���(#�ޞɐ�4�?0�e����$��ָd, P�xy�iw�(�=���J�ը�x�S���4v��Q�u��XI�$�'�������I�ڥ�0]"��ѾZ�%B�(���	��j�b½�o������{H|QI?��iq�
��IY���<h�b�M�e��	2Ys���p���l����	R�K?���p0I�+H�^�l���;M�`�Xsy�u*Q�R�b��DS@������M���gR��"�	\�z�;a~7l���v�G��B��}�N�X�N�#��O��u�Emkyb%��?�T>G��|X�����8}��Ǧ��Rb���ߵdȣY���,(���3��e)~�o6d��R��ް;���ZG:O�4s��C�͙>��>����#ny�Ul{���eQ�e� ō�����0|)�G]l������u^��xLq�2��Y���D^x��#���?dWeƇL9+$qSf�v-�"����q�K�۪�F��N!G�eJb��w�y�g��eڒTzB�����Vl�(vV�h�=ltj�rLx�Sy�ˠ`�&�W7N��7����u<����E7eW�L�x��Kx-�ʭ����5ݩ�Z��q_�wͬ/��Y{��W�^W�����G�o�*nq�;��
�L�4�iSîZp�CW#+Rq$�36��bd��Pt>rޡ�7�4�������amx�\�G+�i�����
5��^��p&~w�D���EuQn 9��4֯L��H�[R�(E�5������L��ň�l 3$6�"�lm���#(����*]�X��85�(�R�,%������)�����7��KL�5_ZT�:�UfS��Y 8���jLWu�myoo���y^���a+��ш�U��-z ������!�)�:�
c������#|F�jִ�(����ېy=��ޠ�����J������%��O|~~u�^&#�5w�;�E�h���������K��У��y�2�Ի�~�Z���S����K˸����\���j�}��?���e�U�M?�M�����i.(�I��W�w�}�
��U�WhtòY�J���֚�ٽ|��Ȗ=̔yW+�L-XjqGŦ__���rB��hר)�Q]xi��UH���*��g�{���u_*` ԉ�&� 9o������U��.\r���'����W��� �]��X�cy%�(｣bJ�@GB�1��[�7: �#Zc?8�+��۹����^%��c$D����* ʗ��C#�,o�,�D4h
���l����7���t����E��{סj�c60�6�a�� ��+����m�%�����5~M�4�6t��G�P�S�q�D����-�������G���z~5w�]L�q�"ӦGS���ă�J��,xJ�+�kl�,R$�v�aJ�<�@��m��`Q,6ۑHC����95َ=i�A�˶��a&�]K�����%@�ᆠ�1j8>:��7P��:�L�SFo[	�%z��נ�t�^7y��?��M�Kꄂ��Y�� u�U����Ќ,U�h��F�}�������_Gj���߉H������2A�/���'&�O�wH�;����#Z�E���BT���'� c0���l �jo*w��ƫ���ķ��e|�U/��}>�S�x�F{�넩����y��5�:��ť�q�_�y^B&��h2+0l�{&�j���̬O����:	鼑$bhX�\͵�(# tg#�ZK[-�r�@_HŚ[�s	-����<N�덒��Ƣ��vÿ��aKq���^��T�l(�qfՒ�}+�<�|.<��h^�30A���%U����WA�(IX2�Xພ�[C_t�fk��숞�
#db��X*�zޣ�ٸ51_��S��'"�؍��72(��'��`�0b���N�U��$T��T���z�%} ���y��|�΋wz����*
�<-�B����g�m��тȃ"5 �'R�90�o�r	4���XxC�nӂ#�3>]~�UeQ*����'�u�RA���1�A�ٗ�i�z��4�r�S�l������U�]OZ�H0ԍ�l)
�����|*BJ�g����<1����	�5iY����g��Pr�,�ϸ�H��J����g-�Ed��J-�
�{u�-gV۝���c���`)�m��9/ǾR����N'z!����n�ex��!�VxR��{Z%x|�J��q�7h"��(�2	Ib�ǿ�k�������Ы�=LE'M��XL�L\�>p.�_��vO�iU?�{'�=/^2�0�b�a�9X"`T7�\���������/\��m�L_����3
��N>A��(�O�3)/i�����e�v5��Ԕ��x�Oȣ�m��6,z�?��D��0����>5��K��Z��$����=HAHU������x�Z5D��dl������145$0n�<�|�'*Q!���i�`P�e+��e�\�[��t"c�C�,�1 �J�y��g���1��?ms[6�����<��F��&�h&xV�!f�Z�c��E�,��R��L�0�',��-���5W�q2�>��6/�wG�:�]Fi��okm�M�^Q�%#0!����Q��"`����ZJJ?�U��Kf�$���LyL�{�=Y���l�2���K�!롚���B,�׽o��J����@�l�~� �7֨�. ��7��&e��VX�mɖ���� ?%kR�� * 7�M�=�Zz���$�	M�MW�!f%;a�卥)W��߷�tH���^�p��D~� ���V�)KM<G�3 N F��Hpv��ջ�=7Q1�|{Ж�~3
�^��7�*�E��>��A&�B�N�>���c�������0�R�~[Y�s��Y_Kt<�U������%��3�FhF#�x������"��� џ�~��Wuǫ�	�)��~X��i��B���Ҟ��?�Aᇪ�A���ò��6y��E&2|/ߠ��K���\�D?R���b��öC^�e)9��8�ـ���������/���Vl�zus�D�j\NW�Yzl]�G�ě+,M��e�ǫG�(����rUKJ�?�B����R^"��y:���<��WA~?s>����Q�G��Ǘ�|�c ���l�yr��e�X��tX\��?n|�4��dԲ�"X���25��JL�=��`Pz	j��ׅ׈C���n�kV�A_�X�f��yƨ󲑎X�r`��|#�A�ww�������|U��ޟ�}dI
̦�������m�����?�+�J���E�4&�?��'t�fM����w� �eݗ�<�՗36��E��א)�"�^&l�M+��ɒ�q��M]�v_�ʍs�/$ɒ�WU�?t�Ձ�4��[jo+#*��T����N�4�4j����p&B�&�KpI��O��Ԩ�棱�̅5|]��ឭT\Bt�w�L�ً8�v�)PB��7��BD��r�}r�OD�_��M^�߁���|[<��b牱�fk~�����7�}�,]6oL,�V��b6x)c���BL��d�K��>2�=oik�5c�-��7b��
z�L/�7��߼�Z/y�ׁ�M�l�.|n�Ԙ��8O���]l�L(5-����a���2���^:5��R٪�P>%���F�v-�:��b�"��O�H(F�C��̮�$��l����.�}	9=VvP5�8��S�jkTrw�n��1�q}Qo3�v?.UIc9�n�6��Է��f�b��_it��-�6�~���ި���;Ls�V	���_zݹ�G��Q����k:�h����Pz��H:'�|^���^!֕��W�fݲ���tiߋx����h��o�m�, �b2������q�+WH�ބ;̴�����B��	�����=�j�%���7^� X�QY�3�nI֘�|Ǟn� �;��7� a�Ւ��c�e�x,�d!H��}G��ҕ,��
�Yn�-7��_q�$�*��0|'�t-����/�;	M2o'�λQۗ28�C�29�|]~U�k�٩2���5e�ޏ�bp�!��@rI�����w�g�ɻD�G������[�G���y�:8�8w0�B1�M#��d�P7�9��?��Vqp54�Çԫ�� ���;\��7�����J�bl����R��l�'�rӚ�١u�Mi�4�;-�ͱ<��;�E�������Kh�L��kXf�i}����
���.�?hC���u�y�e�Գۤ)�f��Mz�\��O�v�	d*T|x��q�)M�[�ԭ2\d�ް�o�T�Q�8]�����`DƎy��P\H�-�g�9
yR�WFG=�'�S]�@��}<��;{�HZ�0��}3�Eb����H֘�OBf��?�`�减@��M!IL�!�P/�e��Q�tf�L��s;�s�8�=KF+$}2��0�NR��`��bu3�퍛N����A���L��U�8��=����%�������Pӱa(j�"����E@2���/'�:� o�,=�x�&>e���Na���'w�u������s�v��d���w}�O!hR �>H�c4�vT��
�L	Pu��I(��� �;�Z�Jx�&V(�ԚM��x��L ������g�Ҋ�>����
�"LR����`:G%?02s��̑V�7=0����C2$���~�C���:��gcv���،�f��-6#�d?������g�x��������Z����>�MrN���".f��Dˍ��9�M`��`�Hd|Ia-�a���[��T�7]�1+8�!@ᰲ;���iyL�Ú�m��'d:�֑���$�3��r�;��~���qr-�h�t_t$�J䓕 �����<���!���X��P�%/R���u,P���DKl���\SeVތ��|N���G�!��C�ں�%y)�nN�uz����[�dC��v�s
g����ª�m��4��1��(R�Sa�j����jGFJ	���}��z��oi��ߩ�Aղ��n�ѭ�IY��~�±� 6?���a���Z� �28d�+6+7�v�&qYR�v�ֿR��o�DI���~&{������ |ȵ<�O2?2U}K؀��%3�\V4S�t�����)l�� ⚎B9�|���_#b��(�<ѷ��0WW)c|��hVq�|������H>�\	rl
~�����o��P��3�x�= �_t4r�7lv���ݱ_F�q�]HQ�o=�G��̰�{�Q,��kzJ_�@��f���Q�����o���6� Ed���gR�Z�¾��7���;��.�``������=ٍkSpZ��u�h��C�5��8�d_lnt_���mO�D�_��s���KpQ�"�J'1�*TQI\/=���[��ޣ �?�/���o<�*>�ѳL����El���#�؉q�6��O��k����lA�)��2XC$�9�+J�I&�����5�t��\�>�S��݊`�9p���%����G����z*��2��ݸ(�s����:�J���O�^��&T|ҳ����]�C�TPmI����ؿ�
p���n�sf;:�l������2N72ǖcT�6�y~Iz.}�.��i�G�[d�JF"�s���j%�iA�Qiȋw�	��& �^�����N���f]�$��Ѣ����p��_��U�>�mMэ�\���Bqc2r���R���dd{7��Ri���gь1�2	�4����o�؅C��]����Mɠ�G`4"fñrY����U�d���B`�`���<�No���NT�\Jc �KOH	��̛6�n��U���I��8�4⬷�� ���x;h��ADS[��i�}�Sv.���W�R�qA
�b��!�T.�\9����"�:�/���`������$�٧pNa6�' �M��Stw�(q%�����{�KG�q�);O1+T�T�ŠB��ݬ]�1~���i�{���d�����y��˪�I��ZQ=���?v�}�qR�!��Ͽx�<��)uhFda-Ӕ��@F�I���i��/�����a�ByI5(�,5_ȣ�ͥЛa����p+9��LR���QG���Q�,����M��N\����H6{d$�V7�4����������O0@ܮ� �ܐ�h�`ݢIe����8y��o��!@jR�o'��rb�
R�Zg\�#^/��������S�!��؛��ɒ8!Z��ɥW��+�=�Bod��� +�c8��Yh �pp?Cˎ_��Dޯ����2���-�1�dal����\�\,���w31�u?h�[Fo�w�m��=y����$���.ENv��D�t�ݒk�	��jCG�� �~﵋���ۮ�/��<pc��u�RO���2��z%�3�}�@��.o��K����f>=@W�[-���J�H��jw�^т����\'y�_}�;Dg�VXA�1J$*9'�^���\G{Ý�H��>8�N������A.{��]>oUҭЃ>�4�B�\�	7�x��R��P��Nt�����~�E���B��R���6{�͝��[����l-����o�7���ox�Qw�퉃�K�F\	U-/cvl�uD��Mبr�R}"�xC�<xj)R�E�G,{�q�^-��,k��J݄��2�}C� IX�#��@@���:^��	!'���$�.�m�����0n�'Qu9����d;�����;���C��
lM(
"\~�����aO�����M�GJӥIY�gW7�A�%?��N�`�=]+�
A�@����X���n�I(y�����:�Z��yb����pK�'ĭf~�l^r�\q���V����R RY��g�ԅ..fvD��t�w5��Z���v$�DeDhZ�x�K�,��ϓ
;� ����I�\�q��0DK���E�8#��/Q����U�B����52�ۓ5�_׵���@L]X��=�;gB>�q�A�p�މ��mCU��.�簰M�El�����;M�x���8�-�_si�h���xb/�-M��Tzs�6\�~aWKg�1����$ �U��?��Vũpy�]O�7ssT������86�CP"�	3iS+�n.���&�Y�L'� �p�c�D��x9�au��Rx<͗N��3�2�����M������
˴���3�RX����~3�����������Ș'�MC�!��2�Kеؙ�n:A�o�0���K٤��%vRw�I7�׶�f�pk�S�ơ��X4/.�<&>��<��{�ޓ=�c�����>���_��V��ʑ��v�ӳ��4���rePۺ�g�wwt��������U���e���z4�x�g�H�3��o�����N=UI����k�(@���Ns�ח��c����5�#����?VB�t~!~���
�R1����_��1:��x+r'F�t���p��7��uJ����1!��ޚ�3ǂ�WJ�Q�5F&P��/5�A�r�E���3����g��� �E�������p��ک�"���C z�0g;-O�NF�b����B�2�Z�-���>�k�D�+Vx/���YX���7�����1O˓	7UP�T�+���i�,�@k���e�-]���(��I�`��a�B�r�rd�g�Z��TC*�o��P�L�������j`�Ԉ1B%��hu��)����_�*x��r'�8$��4��A�lay��RӦG;#TW:��+�dWo��a��݄�V�����]7ܦ��ڭ���s,,��gHi�X��= Ļ0g�6���6Ƞ|���Ʒ���0�xIJ����V�(	�����[oW�~��K��-X�R�v�Q��@��Ϥ���������p�"�5Q����*䥣T�b|Y,�Hh-�)���0��(3��\���]���>��FA�����q'���Ô�ʦ~�WH���T�>3���:�k&?�O���ď@�\�e:���{)���18h�Y�۷�����'�����O��TH�޾�mϰ��_���^;���ҫ�^Yǜ6��UHX�K6WE.�#�s�~��D'����z̋�:�L+iB4|g�S���.ɽ/�ƌ"���:�z�ū��`{���`,6�d�"U��ŭ���r6^=ђ�ql�:���6�0��M�zŖ��N����E�L���N��r#/�#��%�ݡ]%�۟�؁��@g'��2��yz��	L,uAC�h�;f������O���vx, �\�CE2��:V %�gb�S���ь���B�֢� ��)|�#/p�@�oNͺ����?J�������u�"Xz4Y�`���Ŏ��?6���]<}�8w�<���N#O�\�Ę|��N#�@��9͝;kE�6���v�TP�>�Msׇ���X�k1��Z�)i7�$���5o��^'��ē����76��s�}dT�w�۲� ��_c��ƽ�¦|p�P�?Db���4}[�ك�n뭊�(*�Js��J�S�d�N�ɏav6�ʿ����8�s6��^7tp��x�F��Q���b{�$�k��[�Lt55��2�)�2hz΋��hOw��Vv	��HY�e�Ag���;�z�u����eIj ;Zǜܟ��s)�7���H�%�̜4�����4F\����S��Zg�̀�M�KN�#��ˏ�/$�S�9�]�P_n��������R�4!�2!�`���Flڧ7�~z$5��	n�4�'/+�q[�����:7��Ļ�ߜ�΢ʳm����J�ި �`	����� ���4�_Â9�HBbqxf{L��Q������Tq��3<�6% �ELB|�x��@���2r1"��D�	n���U�����^c�0����bJ\X;���e2P�Ȥ<F��&�X�3�w�{�m/.�k�pH���D�iRV�@���@8����ڃ3�7�)�@�eԹ�@�����#6���?P=z�٭����[�8�v�mU��)��ڦ�^��,�q������o���.��ӟB�*^�=��;GB���P�40���x�/b��v��K8TqC�a�.�l=}�nBLx��k��tɴp�Q|�48
r�����J���<"��O_IM,�h��:;s�7h�9���$%��?��0f�M~t;��(�Kcۇ/K"nݟ��	�p�w��]7�s_+4��D3����5[�A/���LΏ������f:x�{���/=e�a�[31�B������5rٌQ�k�{F���0���ܣ�x��
��������dɐ�I�x����������b3����*ً�yX���p�D�_&Q�&t#�~b�èU5��v�B��}v� jf�/�TI)��R�ƪ��m!*�w�!�[�������nu�%�~���ӥ|�o	��]1��>n1��Q?X+�N"��ءM5
'��K�@'���H�(Te�AF.��>��/ox�6�
\S�3Dmmi��J�D`���)��l����{���Xcz��F��|U.݈?:�9�&�>�~/1
��s���,�G�D~bô	ЁbCC��~>�V��h���Y�Qk��h���O��$Yt�"F�r��ƁJ!>�p��D��5�+w��NY@i�e&��kia+
O^U�M���:����;~l���=e�vf�.�"�Go��P~�D� {�Ms�^��9��Hr�p�-��������(�i��2�X�� ���(DP9:ێ��(ȅIaI[;!��u.�4��p�����rK���$Q�07���[I�k�-=ή%����e�������� r����ۺY��Yr���y�Z�J�G��]���E��XQ�3ሊ���cE=`S雴�t��C����l��;=Tt)��(D
��n�E�u�h�}�*DP�鏩�Z�}?Ym�@!Q�D�%f�J{��7އ[�����Ě���F�?��p��2�)��:��I��l��]�ۖp���a,���T�e��96��̸\n�|�}���w���GӤ� ɟ�.�x�#���"����v��'��X"�ou�)K�9�-#�G�[����Y����ZQ��莁f�0sXDz���#m4y�Im�R�CL�΍=�uV���c�o\�ɏx�����㒰���L��s���4�}(!�Q�~p�\zo�t���6�u!��O�A����x���k���WA�|��gqvT�E|�D��9����#UBS�Ț:���|�"�\v�����~�6}�_7��CQ��?0��ڗ��bI�U�!�]ʲi�$�V.SSCӧ�l�@�Em���|оiv>m���>_5d�ZQ(Kzv�V�q]:3]S݁�v:G��j�"ɬ�gdZ�L�G����-�Ѵ�&��� ����2key�ϟu^��E�1�8��_$�A����M�D<p,�p!��avfY؃Y�j/�#	L'6 j0n���p�y���D����F����)cƤ�93�SϘl���{5y���-Y���.b)LH#��j����9�e�@�tݥ�	�h�%���5 B�.s:�s����ZО`�{�s۪	���Ө"ʣ����|��2���E��
O���7m..ˍЎ������K�����`���l��=�톘���μ/�������Vi�Qt�����J�%��ފ���~&�ɬ��>IeJM�Y~).qi�-��4>�TJY��ڿ�2|�⫘&w��6�{��x�{�i���E<w>f�
�@}F��b:��<��vv�^�ub{�,�F��G7��w�K$~9AŊ������V����r�=��Ab�4^R��]�Y�C�滦O5�Iɐ�0�&��|�{7�U�);|Z]�X�?�w��o,�ӎ���	��QV��X����<-�X$�����*�
l��]Hŕ[�e/�ؗ�{�m�i�����<�c(UD��b !3`���XT!(2�&�a~?��>�����/�Nr��3ۤ�v�
��ܵ��=6Տ�f��I B�� [�,;�[i����n*��\�Aŝ{C� 9�4S��x�)��,n�j}���r^Q��
�>���\�g�	�x�����s���!���T�q!�<��Q!�����jo�e	=&_�E�ޓ���i���y�H�c�/����D^`���`�����<�w��Wn{Qo��}��{�)�a}	�d��}>���a�>n���,v�d�Md:sb�ا	<��W\��;��Rz<�u���b=ܐ@�a�ޝ�z0���5�,)ӹ].R�����Q����Z��
3��P��o�b�}�#t�4��3i9���V�v-�tn-��N�
��c �&t5y㛄�E�~%�`�G��t��a�v�.���1eUٺ��[��I�uG%�j�^h7��m�L��c�=LF8��zIe��������_��c�t�����8�*u��������v�y��L��X,�K����5�G��e�i�|֭�"B��^�}XU���s7?ۑ�D��2̣>�̓��ж����
�)�F�b�7Z�Jw7%-?�G�a��a�5�j��U�%0;(I�R�ŭ���{bIB�d�pue�S����c�a�=J]�(^⃖���Ù�����b�b
���\� �[�Up�y�4`C;;���%��q���~��- ��P�ʖ�P�E����B4�5�^!���o���G��j)VOɟ|R*7G����&�%�
��K��V�>��qyːP�i���۲I�8V%4铜g�&�a���q�v�����_jP�.z��j�F^WU0�n~Z��=6����s��c�^�����9��&�ƂQ-�RO�Y/��rT&�u��]8NY�=��O#����T�o ��H0��b=+��Ղˤ������S��mG��a�дM�kCt1 ��H�P��'/���@�p��.�t�%F�D���4h�vN��-S��q=�lz�_�of�����_OK|�A��B@ �u��x�$��pGKUA��W@�h/[��O����|k��v���'�@+�=�����?�'�u��¤��xq�t��_�T>�+9��i�hѯ&t>N �1���(��# 8��%�YK'�sL#���ɛ�dÎ���,�$(]-�L�N���P��c�O�6ּ��/о��~x��B�e��0��rs.�K}������u ��<�6�0x$" �a�~�M��{A��EL��s�����>HMW��w�]�������F��=T�1�:�v�V  ��!&D���گJ��B=)6�]Sw�7��Vh�,�[�ߋ�����$�<��<4h��<$ļ)�r��h�U�Y�WG%��L7h.l
��\�#�cum�o&wCv���_��k+���GR�g
�t��0�~w%�o�T��dP�B����ݿ��:i�j SI=���a��	���w;`q8:��X64��Ә)З���m�"z�#���\������+�xNں�+	e~Ԣ;tl�ڣ�� ������k*WJ�R�ͣ�;2Q��h��,>���q�0H�뢴�ao'����1'�B]�(���3���	�^T����X�ĳ�/�����׬�O��5&?�f���-������#H>n?NW7�E�܁��_�Mk���(W$�뼾�+4 @6���Щum[:�>�	k��N��|1��\����� �0��u���v�1�Id�Uy�Wo��9��bs��9S�y`"Bj�g[��/�Ȍ���6�-�ֹN�ROHV�mv�E���ד�4�v�ύG�P+/	���:�x+	�8qf���F����+����4�a�Z�X�މ�}3��K6M��)����z$K�F��<�����2��M�G�B��h7�U�1D����􉨀/��kzQS��P~�z��:z4 B�����"����FKv�D
6�8dm��kp<�����H��&�W�C�|2c��<�x8��3�D�!s^��H'J���`0e	�Mk� Qf��D֠���>������09��٦����Y�j]�*�S��S�G0���4��Y�tl������2AmV������[S,D�G�;v��a�>�����F��<���@�������<Z�`��R;s��pY�h��B������PaS.��z��DT���}Vo�Ͱ�B#>�_����h���o�վ�8+��X
�|j�
<�	),�.=NȻ���9D�0�V�sVr�R�i�la��ۅja�g�"+`Y=�qR)�?���Jt��>��X�n!bBɈ�T� ���D;v��`���R"���Q@��О�di݌d�Z`���	-��X[KE�x(ؙ��:���oz�K�`3���O���77d�j�l~?K�FwD�-$#��۰u#�T��0 ,8���נ@\��zҳ޴��G�ܻ�&f������o���`�{�i��{�~��Sz�/�y0�t�v�*����N]6�'�d&
m���5�ƴ�@������$��pu�܍�1�ݡdb�س����y�k���`����K)O������;Q/� ��h��?!��]��٭�p�	��a��O67�;Pd���ց`�7�Jc�<C@��L�& ��� ��Y��0{[�q���Y5zd�w��9K~=�BV�q��.�f֘_N�����n��V�bݦ���V��f�(f|������?{��1���ڝ��́�wD/NB��fo���JuZ�X� ŚI�x��ކ[R&��M7.��S�
&P���߿
c�]dڇ(@�YR+P�[YX3�u]/t:�8u#�&B~�6�!gSa	V�����T}�~Jѡ`������o��7�P��{�)m�J���0݆&o�F���!�P�3�!���7�IU�d �	�P���q5��U��K��6�7J�l��e�	bE�@����'J��8
i=9�v��^5m����~�{�6��Z ~�a܀������#�����J�+�.�j,5l�aO>Ř�����P��45��t��R� ���a�F2"������1ҙ���L��gX�(Ω�U����2;g��I!B[2i j�(/j���t�r�[PJ��Fzty�>��zu���,U(�q��]lѦ)�i����.��������T���³��5������2�-���Vçy����L�hE|d�`����P��HW��¢��N�$�)���C�/���(@d�������G]fSs�m���i��<�9�	-���Yc`#\�zE������%2%�$z��^��g��������pܢ ތZ��J8�ӵu��r�Y|�S3.���q�W�S�59E~-����[P~ցqn�������ܫ�G3=L�⓲���=��v���ΪG���`���ȝX��.���Z�&-��)��]�;�AZ��j�$����$�\��!K�T�k�st�犁�r���>��w��h_���ÒG���oO��T\d`�|wۖ�r�ԟ=nN��
����it&] 5���f�
Q�@����5�9O$��$?+�z��g�h zgMʸj�ؤQZ�s���aR�O���mDw%c��7*��ՁB��c�{,��L���^>��m�E��V^�5�a��N���@��X������.b�)iٓ"b��˼ġU6j/�6J;���mP�ɯ���tQ�BVĄ�bN�۪�����$əA���fޜ@+y��$��J"��ĝC�.��Ե�gJn��(P�5+�/?kb�;��32�l�п9�:��@t���U2)x�q0�[X}�|�a_g&e!?aK3+�A�K�3��BN��^�$x�+?�����&W��𥅯'K��_D8�d/�h�6�>B`�Y$Aۍ�����nI4Xɓ2t	�{�3	χ�+�q��t&ʘ�փn��� K�HU��﬏lK	<qI�AZ/Y��_�f�����
���D(qTT/3(���n�|�yӎ�:��gW*)��l"`"'5�����&w6a�ȥ�{���k�mwBV��^�ǂ�]n�!(�$��qɆS�"�M��xٹ��|!�V/ ����zkZh�i�)ᬆ�=7�";����\bl*k��R�p�,��7�����i�TE'�3r^9��Z�j�8� ΅�"6�/m_��V2�B(#͢�?dl<�3�w�6�ԕ�nP�0b�h�Z:���Cĸi? e����O������B:�@�I�&:����_1�;L��7!�n�鶊t�/vX<	�2ktD�' K!��":L�ֽ�*�UDL�<#����]&,<�N�A������U7﫨3 �M\�L~<�{��v`�f���zGQ .�NT��/��z+���#s�x#��C'����������DiW��V��yGi�C_Q��R�vi��x'�MQ�w�;����ɰZ9�I-�C�#K]�R�	��0����7���-���+�*Z����+��㏉���4wI:tL2�<��$��ة4��1�0���s����<�7$ʨ�_p���@�́:�mn�οqȵ���3Юn-��a�Q�H��۱Pռ��Ӿ�5Vɡ��X�����n4+�1c��V*�C��-��5?&@���"O�;�:��D鹉���"_����h���}')D-P��V֟��Ί/�V#Y���]R�'�Ӈf�i� �n�X�g�u�_��aR���i��O3���l^6A��i��������U�^�d���+ޗC��K\��N�J����J��Zd���±�� ��[ܨHY�[Ηy�G�T���]_1����)���{�@��q���P��̜��V�����K�C�K��@f~m��lygA;��ŪX���<_�ո��a�9�Q�*V<��r�29�/�O<�0�����	����WV�혠�Y��1EWY�(������ψ�r���7(��� �u�X��a��=Z/JݔA3��$e�9�9cs_�
)�K1�Qw�q�eb�@����7$�W��
�}��ɻF�X�3�������y�����e�3�&������4Iα�GUs";ȓ�MmTO�0'�3Ԩ�e��P6(3I�a3�<8'�
��m��()|k����k�-Ⓢi��|n(�d�	(u�g�������K�at��m%�m\�<��4Ԣ�H�D��8 �<�N�vl=R5�=����kJu�w�#?U3'jdS�=0��8�_��
�=V�j�7��5��$��oeT�8 i�`��]!?iyڷ�u��!:��k��aOFP��,�����0��s�l=o�n��i�L�	Г�H�>`ǥ��8A
��Y��,)V����A*f8��%����V����5R/�+�ȳ\�TGd�`���*�p$N�*`�c��F��2�eS����� ^�ъ��j�w&��ם4LR!`4�O�6�˰7���"C��v�[ D`��.��r�յ6��5���DQk������x��oN��<HD��8�BU��}��7g&M)4�MӵR	HE�$ؿ��u�W����@�z ��h"�$V���E�۸>�i������|�yl�y�Z���갢{��9_���P�K-1���$�Vu�|�~=^���%���Kh�
��ׁ)�jϮ���( �d>HsS��\��ZӰ6ì�H�	� ��|c�d���V��lo�!5.��ϴ���Hw-�+��#�����ί���T�&I1��������'j�a�׫�w@1qCBb���<�Q!��*e��*��?���WZ�)'B��l�1+{����7	�R��5�fV�@����-��@%Q7����$?�ZM^�M`���ʺMތ/�)b�]i�X_t���讣]�-+�L^F�ܤA����xɲ���7͍�	���5������~[��]�:��߈»�ɿ�����/f��ⶎۀh��8'e��Jc�&�l�/S��
h���R^3̤�w�[��(*;��D=����`:����0�������O�N��-�q��W����^�i��1�V9��c�1s>8�9���R�~Y���d,�|���ƍ��`�P탻�����r���P�8�g���c�};�;=�f�?[}�U˛]���գ>�������tHl��g�X�'6�GO�` ���T�-��|�5it�
�e'9[�E�jg�~ܳk�#�_�}(�Q����\B�6�w�/�>#��ߕM0�ܟ�At��2�f���Ϣ��d�Γ9��=�����X�?DP�@H�#O+�.m�x}$j6��:�5Jm$���D�ߌkݓ5b�L���������J�D��~6��y���eW��7eCN.F�B�+CR
��}��~S�U���PG�O�e�)&��K�������J�Q�wI���õ�I����Cįk��������}ٿ�u��X�a/�9�dgO�G7f���S���~]��mѓ��&16�5s�5	d��_K�UeM���{Q!7���'���B��2��6���T����;q�
���2���Z�1�~ �.-�01@q�G��n��CF��f,����R�����e�:d��PC�c=2�u����������~�7�Y�/G��\�O�b��N�:yUgF@:}�<�\!��ٶ�]ا���%��|nJ������\�z{��s��(~ U}�G_
�ܾ�-L����5)@㫪4+4�гj+��k�l�o��-��7���櫩?�Oi>���;-�<!�W��b[i���0��Q�\�>�س��c/~0�v��}<������9�u�1�2�1v!F9=�>8#y"\��O�@
��2�x����X�&�(}�"�B��(�e�;Lk�@l�Lk�c�P���(_������u�y%a@��G.Nu��&f��cAM��.��HF	�T
N��c�������hd����+�+�Ĳ�W��i�)Sfx��ow֛B)��SK�e\/�]����jdͿ 4o�z��;h�@�:c[Xp*¥Ӻ�2����§S�Y���*`"�t����m�'ɴ�;u�9��H�%����)>�0sv��Bb������+�%b3�ɠogB����n���?%=�P��z��NFY�'HCW�-�p�&p�V��t3~nK1�����q�40Ln$��i�ѷ��>����^�Ne��A"	�d����<��3�H�����ͫ7v�	U�J����,��� �A�����V�_iwѾ9�rI��z�+W=����n�ҡ�����.pb���2�R(�<��ug%�������篤��',)�y�]P�����u��1M�^�G�B�	��{%l9�xm�:��N�z��f����ܚ���>O� XquF���s+%rlQ��I��I�&���-��̨j�9EcD�y�M)`Y�a��5*��)+O�"X�.^�ES>f��v��=��)�"W��dQF�J$�!�-8�����̴M5�M�xJd���ik�- �A��Cd���55�	C؆Hr���зw��� n_�\�J�NQa�d(#�L5���;�x�U�����gn�a��%D�Q	��Ҁǝ�E�E�H5@�K$ې��r�FG����M��Ym�.c���@Qӳg�P8�RuY&�(;b��Y'�jX��߹��l���A��ci&u��G���ux[u�G�S�q�mؚ����|QT<M�Շ���Iy�"#��e� ��#�#� �}F��a>j�=wm���V��E���20����%,��q[fn)}�jZ�F�3\�j�a{�1o���g0r����3bM@�&2 m^	�ɓ�?(��O�b�-S�˶�!%��\#"=�-Z�N6�=�V��aPi�;Y[#��ȓ.�ޠ���L��T��s�w�f��b^��<�lN��<��l��8hNB�Х�F�8,�╾�'�x`
�;\qd\���K�-'���L�w0Û	��N�jTX:nd�y%3ޤ�`o����/~	��Smp>Afw�G�K]�$H	���-�<�8&bS������}�Ѯ�'����"�@����o(��ys�������cWm6@$%ͦ�.l������ӉD#qI��ó��Z��ҩS_�􊜓�K*l*�a^P�5������S�����MU�ӮฮPS`�j-��c+q�q�V�#N��(J��#��8/�H�v��'��B�x0گS�(��n���y!}�ָ�v4�_j�m�Ja�r5Z��� x=�^"�㮇LE �s�alb�$H�YԜi�X�Wު��*m��"'U"��أ^��l��#e6wB#�d��02�|�����%��˿JjȰw�����u�QI���a�����c3�-�1v_�\�#=ԫ��:�q�� p���Ac���l����%vx^)��l��v�8�l5���&���H�f��G4-;�i/?�<�S������p U/�-S���6j,vw���N>�]L&h�#�DtZvf�A�w��A�d?F&���!zc�P��+���3V��_��8���6GdJ��ݾ��P��q��2[��������@���0}��H�[�bO�z���u���h�J��<�]qP����"1?�!E�eI;MdHO
s5	���ܧ�>��c^�>��Ֆ���]���x�� `o:3��?�}��_m9� �����ahmݸ����D���]�@��ֈ������s�|!U��-$�X�������O�G���ğ>�J�G���}�����S�?3����>��gf�3�l�5��{�Pɚb���1���v���&������e���!E���␞�?��Wk��l0��㩀x���ƿ2By�1!�1��1cp�i.o�DϧNcwboQC����ׇ�X���|fe�����5��Q4em��»�G �UJ��Q��C��mЋRS��&804f�g��dq3��/���
\�}�i{�Pӌ�t��we��!tܲ.�SRኋ�d7yb(�+�͆7S�? �}���3Hƛ�!���+u�P$<̻�sc�����S��T�5��kE�[n�e���qy��6	�K���E��Ub�!�ʏ4���2�38�Ng�s�!��RS-]�K"���M,V?���-d�t�t$�ԿNW��I�R��o���t�>*�?���FtZ�t<�q�2�8(�#A���
 �N�]U��WՓ����/A��4�3פ��Ӝ��!`@��s~��Q��X_�]];���q�h�B�v�����5 ���$��ayV����fX�&s��)�
�M�.V>��H����ʵ��{K*�4�J��CԶ�א=��\J���s,���6������lE���ݐ �%�w�gVd�1�A�������g5{_�m��F�V�����]�`�P���V���(#�5��hp�bc����B���2�8����8m.�3[�Rapk��6�J��b-9z�n��z�,��.�Bq�&E~���t˽)lR���5�N[��%Y�l�!�|z^̜m[;�g�a֑	(B�-b��m�[-#���˩Q)��4�ũg�t�����F,		�x�o��9z2��|4�x{V�wA+-]���R��֒�Z��ҥe�tV����\q4B�������N̓9 ��IǄ��"w�L�~ ���mȕ��$6(/$��%Z���S� =3��w�K�a��3�V����u,�>y��aV(�_	�x=����C���ql��"��i�u-i�C�.�іע��c��W�z�=�,;���0,�~e��l�WqV�+>�!��#�ibm �Ờ:&�W,7T�>+m����ҽ8nѳ�B�$�ڥƻU�I��a�NB��	����m�b��E ��=[�9����������ơ��1��۴Y��9�>au93� 	RތX�ELE��4��ȕrѸ5��P-�x]���e�&͂����K�*7����}���.Z�j|���c\=l��^u� ���+Љ��bG}&����/诸�T��03�Ԣҝ�ۤ���aCW-Y�ʨD��o-@^�Խ�a��8��T��&���2k��n�Ѐl�=i�j3�tL㪕~"2�k�v�I)�'K6�����kDKy�����a�͊v�W��5��2�;�m�Smmʌ�@lñ�F�J���D���A� I9Vq�����.���$��.�L9�#���_�sH�(�p��8�8i��g�ª�o�f�X&�KγR��=~F=�a6��F��C�H%K'���ٮ�vF���y�+�L<V�_����:N��� (��S,��d`Y��L�`�>^���Ͱ%��H�K��t���ZE�Hw�{�<g�q���"���m��>a��}r�š�(}t�!F"\��L+��tI+.���z*r�!���/u�0g���2����p��	�������%��d ��v6�����E�`$�|W� U�CU��ᑸ�
j�J�AM���h���/�|��S�L�_3~��\�s��i�@�$4�G϶��7M,�Ei�5'nQ��Mbb�Z�ɕ(3h�pr��|Nd�(Wis��C��� Z�x�Z���C1?sT��c�)�D�&Mp`���'�X{d����eb���v�E�s�H���s%�Ѧ��P�"{Ix����@���sI���@|19�srs���*� ræ�u�g����,Yd���p�'�E^;�3���As�R�K09<�*��-N�T$ ��R�y�Z����� ����壢��w.�pL)#)�ɴ$`�\�]�`���-q�vyW{l�"ĠXa��A�2j�u��zX�`���B��Q�	�[���x��r�^�f�Z���L�fr�	��6�|�V���:���K�L��;���F��9>˗��E5b�XO^�I�37�Cv���b�4N�2���N�Pun��c�t��w�5F���9��=$��|F�Ѩ�����"t�y�J~"/��0�O]�G����*��wԵ�@ف��Z58��	�Ȳ���mr��&���,No����`Pe�B�'PU�(��WFl���= 'mu���q��A�:ف���
o��dQ)yy�_���%�H��T����Bg�y-ۙY̝qӵ���,�k[g/s��-X���G�Q�R� O[�1�g�8r�u�����[%��Y����;�]˫��.8,�^A O���oi�B������u�/r�=�8�a�g6(G9۠B�5v����,����{����
c�Fp)?{Q�\#�3�Wg<r����I)��M1���*�PZ��a�.:sm)f��aC�RB<`F��(��
�W 7-�N�ŋ��6�������GK����8�#X�x���h�(Z9�U ߖ��g�
�C�X3A��1.���4��v|,��+��:xޗ$��d�;�p��Ҩ۞�3�&)A� $���N$������]�{Rǝ���,D���5�~r����Ts�����z�����ti�.w��a��O{��ǋ�8{�.�0;XFT�M�u�6䡹+��[�,��U	���iB�@��� ���1�u
��V�H {�6#c�������~���/;�+�_%t󊢷�w��k�FR�^�9�V���ƯjT:��@�0�6�|q
��A4cV���ۄGa����C@vHf�ͫ�����u��{�f������5ڢ�,>t�/��e�]8��ҿ�='ZA�3�D�Bp�c�Nx���Z��{������q�.���D����Jz�8��0��23Y��G��$sH����Ҝ�_����.���!�	�bdJx�M���q�*�dcw����9%^��=
l�Ʈ5LD9���|�\�AkroA\����7�k3z.q�AA�{��RY�����n���ĨHa�ϩ2�����ل� ("m,�^G�
��4��[�BACDN�莸�B�F��9��`���� �����#���i�J�|�wz��z��b��U��/����1��&��shY��b#t1S����@�*fI�|H�n�<JV�XБ!��-���Uy,;\s�6;}V���`O�s���3g���"s*�D��Z\��'��ɝ%1`��Yj�՞�e�y�X}B����_9ƪ �!�X�a`�GC��h~x���g��oP�ӊD@�t���`2�(	:���,i5�e�]�9 kQ�G�h����|��G0���g�r��q�Z��Jy_�oz@�[<9�^�B�L���D�����`��=T�xr,��G���v	(ˣ!�x��3�V~��ԋ�Ր����z�7��;v/�4��U"GV� Mr�����sA/�q�'��')"#S���N���饒
4�E(�4kM�I���u[��I����:�|����)����D�aP�H.$��l�'�+8�K�yz��?}��Ӯ�w+�迗7�����>�b(&}���z,�vv}�f��݁顱�c��𐸯���LZ8�Ŭӳbl��S��W�fO�$N����x������%�
zc�M5�&�Tec�m0%gh��-��*͑gٖ�;�5���$ߢ�[�ć���pg�;��?(����@b�S`	�*�cL�G��6x�Y|	 ��6a;(G2�/�d}5Xb������������o�z[�(�V�h2B��f�����I	/e��6�'�z%S��)���~Π8ً��� �O��O�=�h}�/�Ӏ�"�V"�2�
Ɓʛ��jm������i�V�j�W[6c���DOv{�z��a	cm-�%���TN�%R�H�K��7��L����}���q8��t�|(�4�*٨G1�m3�7j9=
� ����psS��>�"gH>&�Oq�M�)fciLM��;@K,��8��I�^Y��YČ~�d
_ �����c>��n���y|ؒ�h]Ya�{�LL?]�:v����D]�9�]X�Ɗ`�E�J�|��Y�n����ƐD>v�s�� j?{���`��'�F-@�	r�8
�>wV�Z��U;[,J�����1t��N'�Avs˹�0P[&wu�LS#�7��!ѵ�u5���
� �L��@�׆:��$*�]!�Z� Q`�2:�N`���+���`��r�ȶ�,k�����v����-�u�Ǻ���\�[}7WI��r_/fc�x:�tӸ�vMC/E�\1)T��q��
�����u,1:\�M4� !,f�;�yςW��M�+N7�IK�L�\K�$.j��s����n5�{;qt�����[�؎#�r.z�}7��a��W� �'��?���kO՝+�r1n�;Yc%�b�n%��YHU���h��V��-׫-��U����K�Ř��P0C�S8��W ~Ŏ��K�uH��K�5�9!�K��:��;�����tS���Y�]� ��� �i�	�U��`K���͝�-6�#O	�i缚r���y�D5hj�w��
V�4]��Hy�		�������ǖe��Nu9�Ղ hK���s"�l�:z�sq��(o"s9G��nTT[ƮeN����)"ާr�$ህ��+=ӣ�cN.~>��L6[#.��\�$���|��U�Ė��!Z�L'��E�u��� 	�.��; '�:ӏ�P5��fS&b�� �UYF���"�`�!�"]�tz�Ǡ�/�(^()]��_d�|�Wb��Ľ�m~oyJ�����w�>tp�����3�䐥�F�Ͱ�&8,:QQA�0��~?䒧e�P�#u�c�����b����L�\5��b�vːˣ���L#�޴x�5�L��	&Ѩ�Z:�4�@텫����5����S3_��6�A�:<�Me/��$�c���]ͩ+���[�eNÂ�djW�*O�F7��*'D�ӄ\��ಈ�:k���#�a���K=�JB#�z�oD�4� ��\V�TAw���I4TȦ��Ŀ�g��>��LB|� �v��~�!����Ȝs�+&3�j��ħ�v7���^� ���vK�GČ�n%:��;3gX)�Hqё�VJd�#?��B�r�Ve�Z�D*�eCZ$�z |n}rrJ쬬.)�1FO�% V��W	�#7����i����N��6�?I��X;����I���6\޴�1�~��j8é?�">k|Oyzz�̝C��x�}���	�#��{�o>�|�!+yH�?fJqG���J(�Z�H[$,�����*Z+!>ȱw�� �t M��
�Q���#O��ؑD+�{Qz_riq��+�g�ME�o�@*$?k����BJF����`��_���۝���ƞ� &�d�c X�����l�x�Ēp)�"��р+'n��GʽU?	����'=��b���0>;�t$��i�6^S��R,+�=t���Y¸O�f���cn�ԖT�-Bڢ?l����?��M��Bo�+��J���Mq)���j�HB��N�����鿫���/<�^Yh�_��g�&�MQ�h��뽣*�*V?��ehm|o'�ʫ0N϶)�ȳ�0��^����s껶�/R��Ι��5umK7�c%�3�j_���)�'��Kl)z��]h:X�y6_0?$3OyUwa��<Š��b�O�=����lX��މ�֝�z5���#���Fam��԰H����y�t�)@8�!������fB>���~��Z�������\H��5�����c��Sۥ�p�b�}������u>��'v��ڱ`��$�\j�P��@�C�Ҧ<'�x�G B�p�JJ��{N��<0���P��Us�,�^o�.gW R�oJ���%��z���
�h���E8��!uC��G���⤷�։������IQm%�b�w�(�x�,��-�ٍ�$�����xVd~��30�#�&oס�Ćէ�����$�_��j[�d%Zj��>���J�5�ޘ7� �Mnѿ<�<�c`i��śm�(h���X9∸�w���"��-Ϋ�qN)+�qͲ���ٴ�l��D�^����������v�̂�_�/QB/c��[�y�2!�M��5̦B5l�,�W>< l/�n67�H���O@n��i����"�����_���|
6��U�ˬ�e�l�G���E]6V��	"�`����5�RJ���b\ "�&zc�KgN��EG�<U>�}�<u<��[�Ly���Y���r��S�z�vhN�D&fE}�?y�3�e"T�l2�ne!�-��*Lǅ��P[|[���
���O?���L�灕���5;|Ǣct=���/BG�������+N�2]���r��th_�?f�m����}*Ie�ؖ2þ�.t|��T�L�|�!⁤K��_�~3F����{��Ҥa�oDpb���=<���<��ø8�E�7ۅ��M_��=��'G�d�<�:6������*������(��p��E3���K`��fM�|�Y�[�6�7+T\풒R�-3=�������N��u�Zj�D�R�=��ک1|�Ӂ�� �أa���]�^�E�l�eq��o�6-G��r-�m����:&h�O�<�х��M���U��,|:"�`�B#^E�GǓ�B�D����m-FB�|iI�M����`�p	�[�"a��t0S�M3R^�o������,�91+���>AGY�p����yk�I_��B��j�$��P�'M8J��W=�������k@ˆ�d��,����
1���b8>E+Ug��D\�;�Oݰ�)盌�@S��vV�4���i6L��(�1����%W~p�ثǕT�N�I��bj:�sDj�-?��$Q!!}��]'kz�\F��0��v�r+�5�7g�M����u�k�S
������ы�t����u�A�7ԓ��VAB��6h?�ov�Qh��E�꘍'I$���Pv�<t60�����z��'�UE�����L��!��~$��T��nM��}��(��]#D���7��U���J=�O�� �T�'W/i֧v�M�ЩM)�xU߸�bz5.�گ(|Ǩ]�r2eL��z�5Z���0��-��Cr���:�2��jtz�L�e�^t�a3�e�N�y�,{��|����I���i{J:�Yc��f]*�(�n�>y���,UQ[��:?L���%�k�ʷ�]���?>�
���CϤ��b^��%/J��Q��C�G\��LS�\T �t7Cw�4��4��퇶�R�
sPO��Gڎ(�TҁVN����\�\�/��W����r����RT������v;�z18>�΃u�Y�r`z +�����1V�;���6p�����S����Y��~���h���"���Q��U�:K�!�vG�D]��=�^�@lw������F:5Om�8f	?��챌[��!�)�$��̥��k�Ϥ���b�tj���	˾�*��բ�j��8�uq����0K�,9Ь����W��Z��oq9v?
�g��yOCׄʓ{���ęo���;2�S��H�iib�}��{:�d�{D�/�r������g�A�uX����?��tm[��Bn|�\�<��$>U��ۂ�6I �s%��s��K��uwBd	5s�^5VU��l$���l���|,�k�����O�2���y�>���R���k��[�'����J'�@\�{��X�l��N��=d=pc���0o@RI'$XPb�J �CI����/�0f������f¥��El�n�h�AvԒ���N��ݩR�M��=r��a޹h��pA�eOk��X�6��A���Z	̴��-��q����w��nP7��׸�Y�������<���&B��R�f�n}L�n�S��9R|4J��n]Do�1*��E�����#�YO� oܿ��b�4��E%.�� מ|!����d�Wh6���)�i��J���S�?�ْ��%{ݛ�dN��*���lPDmY	���2�)Ԯ�G~݅٠r�t11Ԋ�&��JJ<r ���V1ע���n�0�t]0�}� "��@�`� %�e�n�w]�~KD�E	(*�W&�\`�L�._��&	�`SYVI�4�t�K�A�(>@U�d���"Z�������=GD���S�)�%����J񳂝���w�6D�*'������f�����yC)\SnB��r,b�1�4��5Y~Wf�\2�.f�.]������39�K��]O$)���8�[;{f�?<K�+�v�n䢪�IK'�{V�V�K<�]-��b���j�e��\���O�t�Z��N	"��!�>�I�k&$�����Kb/�.Z���3��
?����sP�B-Ov_!�C-n��6]��hV57��k��l䭏�05�*�T}٭~���>a.q;z�A!�����������x�a0�v�����ph���_�c��W5�7�`C} �x9�w�<� ��C��Մ�0����G�I�9�M�G}�rD������G1�嗣$����	j$*0h�v���'����gh�]��P /o���{G����Ňp�x/���E�i&L�V�,����^���o�:���}���";i�Ʌ�'/hؚ��[���������[U+�)����a�ҽnH����O,��5"j$t%��;&�a���:��Z�+�Y|�XK����Γ���N���h=g泷�S�Ra��D/}�#�鸙�K��Rl��ܣ1�F�O�Ƚۍ7u;"7��2��R�ՠT��^���$Q�z�D�o����64L��>l;t�W�O���AF^U�,&���4[�m\u��#���6�^jx��U$��a��di~��]�$N$��f?d8������:�Fnd��C�]��"���,:��g��1%2���	���$U�A�[L#�#,�{o�T����ޮ��ƞ(��6��X�٣ԡ�zI��m�[�-H���4��V�h1C@��!�|OIƾ�{WU�gz�B ,q6Z�S#/�@P�ٵ�)Հ@������>�AG$�zˊO�g�Uu�I�z����e� ��+ncepYX�!������p�PP!;}&6w6�x�G�5Ϛ��D/I[�(,����[1@��D��{�Q�������Y=�3�-�ߗ��*�Э,]i��KC-9�7�4�N�VϏ0��8�M��r�p��Z��A��Q7�s5Ĕ$,D�?}B�Nwt��G\���֔���?!"w�H#�A�':."��EP
�����KY�q�I�'�l��|�7�1[�wӋ����lI6�=��<[tXɷQ<E�X�gc�!�y��Iaw.�,@'�� 0��r\��-RQ�;�I����(?L�|nP���A�L@?�C����K�f�9A�Ҩ�;ZR�Yњ���������)���W�{�0E�ʋ%��H�
�N(o�՗������!e���m��+����4H�Ǣ��(`8'QmN1[�d� ;�$O�«CPp��D�6{\$W�8�'`F�����>]&��%tJ[�pG��(gLRy'W�0����MPT˺��]e������$7�����h��B$l��`4m��4�f8��w�/9;���Y�ʢ�ZU_��0���U�r�t�ýe{����%kb~t�Ș���v�$�6H�	n�K�+�Ė��B�X$9��<>�M�F����?`OV�?H����=%E�ʦM�MΩLj�����So/w�Y`)~�-�+P��v
5ky>��H?9�tS�0�
n�c���0
��
i�v5�A�S��uL�Eў$~81���ڋ`^K@W�om�0����%/�F�fjN�;ըH��"��H�"=>拝t�_2��C�e�jK�_��������|�"%_\���t�E7��r���6'%h���#g ���J+���������ߩ[~
q�
zDJLH�2�!�՘MYƤd�a�]jQ��z�Z5m�U��]�6R��n���2i�^jD�1�fh�z���6�%��הW�fZ
�߯�.o@�li��h��i�e����u>���v��k/��󋒇��S�C:{E!`��Z���=�o�F����EɿeM�$-5��D��f����M��B>��/BZJP�;M0��RiXa��u x�;zt:p�ͤi����`���[�MV6뚸�-Wҙ��u��!��a�%_<�"?ZGB������*C�N��j�y[�9�1����)1��)!>EWr�O'��ڊ �QOo�5!��f����5�X��𼮃��c�/H.��^��6���'}��j5B�k��q\e݉㊏-7k㪿�:��-ǐ�c�����%��zߪ�B���=�o����}#c �c'��Q�H2�ňK%0��1*����Z]�f�!��aK���P4�@y��p�@��~�𵪰� �JP�I�����D-�ܣ���қ��ىˣ%5�.�����g�G���a����W �w^��<�k"�:�f��u��𭯓\i�oy���cX/���Ǵl�'�j�ߖ����V˿T�@�NGn�1��yd�Ԛz4)�R �T�1�;Q�}����U�=y�]-M#��)�K�O[�r�����he�4:�ѫ�7'��Lޫ�krB��ҵ���O���J�����i�sK�U�$�P�4(���gA����9��1��HK�������;���6�e'dLT4��!l���wW��Y̐���е	x"�4�.r���S�Wc�S�]���F��:��~�1_q7����E�.�݉8�z��^����[� �/q���M�o�6��E�d2'������Δ]�'���)Ρ�C��F��N����۴P2�I��[[����]��r���y����q���̳b�*x
���"��>���#�*� ����}}	A�@�3<�V3K�l*�~�ik(?r��ർ��S���.m����M�w$�Ǫ���Q�
t�o���7�%�=�ڔ�W�9���R+j�yc�/&�1�>���]s���Ͷ��`.	&��,��N6�����`���ۏ��;0rj#�������2K�Me�'�9Ar�sV��o]k[�M9 �+�3+
<�O�IE�f1鄠ۇ;�n�P��+a;j�~�4���n���\�R�s�����2�F5@�ש��M��ڜ8�J��#��}"�8o��Y���D��'8 �� ��*�b'�TH+�n,��h%FB��YI�b�n*�0�A_<�Y7@�T�&�"F/�E7�К�p���#;�������e��HQ�Uh)0-���t�ޓ�h,b����RcI""z�6��P�`l�C��{6��E>��� U*DH�l����H���|}Ǐ���u��QR���*�[?$�އ�-�f�/���1ⷉܼgY��A�{����BlFdM5��/�
���B�&�~~O곲�M_#T�����h�ǣ�GmS	S/��e���&d���=��k�8�6�N���q�u��9���y����@=�J�z>�H�6�m�X}����	�Oh�X��!�X��?J�'@E�4[�bH��jK��C!5��I���_m)��TYǷ�px.�E�|;���6��}}���o<�R���SA:���١���?�C��ӻ�Z��7pt��tyLIغ�Z�����ze�|��*FII椼E`ix܊�2�A^�{��������Ӵ�4�x�m���|j�U��5sCl:n����dm�w�U���,J�������	�ϟ���)'%N� ����ى�D��K	���-�\��X��9�MM�!A���6@s5��j��n�dW��T\/�֔L�S��a -�TP�dQ�_tO-�1.�?E���Tp�Zx�����_��{�g�F��Z���h"����V8�Qq�\��+����p;�,7	ؔ]�;�5>�e��qC�� ��J���;�W�~8�.�?�@n�'�^v�9��=��=5���}��}�ӝ�[6�#��<v�J;&*��x��!�,��F��ˣ����	�<U�=�-�?)d�S7�*XJٷ~���]���;6@���5��R 4I�s��1�r ��Jii�m��J�߆[I�XFbgU���3#�%w/��P#A���[�)�t༯��pD�]ַؒb*՟>�)<�r	�������|z	�\Џ��r���-�����)7b�	Rz
�y��)/�`�֧���#F����`��U8b�Ch�;�ߓxJk�n�8
!�0Q\Ԁ���o�V�ݰ�f�9;R��l����*�L$������'E~�݉,� ��"�L�x���6nxu�L:U����@���I��/`�.3�m9��F�K���֞�h?d7���g��ͧ�Ae�"ߜ���&��}h�t!���9���0�2ϧ��Ի��Z��s���$��-M��ծQr������
��h��r4��:�MbPo��Eb�Q�۹�1�,րǗ��FjT<��_"	:��=5���q�%�1���ޕ`й���+�!��J,��#ls���%Ջ~�}V��
�0q�H��n;q�Q���vKPl+9hc��ɸ��m��rz��[j�.G�vJ�G��O�wd@�uL�c�i��v���#�'�=5����;U��+r{��sf!mv#����9��&/��\!1�`��c+�F�Q� �)�U{�R��|�Ƃ�ʒo�Z�f�N?߀]�z�	���RWR��n�7,	����݀�d�0~�86A��a���2i�%����)]����ré=�~���u��Sa|��@�*�m�cT+E���`z-sO�+�A��)�kym��+&�����t�����C�(��š����
N,p�}a��Q����B�㍼�����P�b��"r�`ݲ�)
F�p>�#��Z��ѩ/42D���X�~E?�P.6���&t� G��=�J�Jm�b��7�۞VBANk��iG��.����8�!�N�[�i{�+-W,^	ϑ`�R��'��J��B~���o�L�����4� .b��c2le������M�d��U��s�����2�m�2�~����;����h��P�8#Pn��󶉅�.{=n7T�ᩆX�uT��2��L�ˤ(���|��H����~a98���炍��R�4÷
��Tl�h,>�^؅�2T#�-YB�9�K�o�=�����1�+�õsB�z��,���[�q��:��T�V�7��[��ȹ#�E�?[�0A�Y^|����ʌ������v]���W�O�#2�gI�Ҁ���+B>
q�*/�V�yP�7�Z>iX߷V�o���&�����UQ�A�����ݲ
k�"�*#��Fh���"�+�QoL����u���D�Y��"⺠�	9��]�X��c�����ܧi	�t�n��,��m��Mn������3�Jz�9���"�_��a\i���.N��̂��e��f"��Ŀ�rx�"]�;�B�N��s
��`�?�]WEܪ�?ӿC�	̞
��D�1i�+�=�(ky4{n�s�XrU��r�)�>����\j��bӯ��a�'�쌐��C�¯��NV���c��2V��>=\O�Q]�ې���C�'5k�Io$�R������^4��ҋy�Z�Z�B6q=���-����R����#��:s���j�6i\���r7�
�9��X`�f6��P]�E�C8j���q��,�N�F�]��������m�(a�>��]��Q~���;	�M�}���*x?�	RBE�8�N�Z-��	�`gL���صLs��
%1��3+��[2	f�b�P��}�@J�d�d)���X�������B!�7���c�T�mI-W���~(����|쁘����Ҹ	 �
p�e�69t��)&��t&"��m�L����������^f��� �DS��"]��T|Vb���<=��}��B�%���fɞf]��K�~+\e^���H��a�!�[���ȍ
1p�ւ�֞�^�H~�Nq|����M>bR7��[��(�N�w.=,��k�~X���;�(mWZ��"�����x%��� �����;L>��x��'&�t�\_�> 8�o@�^ec9�C�?����p�Zi��He���ـ�'�8��K���ƽ&ġPՌI��D�����l|���]ʋ�>�����n@�5��ӝ�۲���3��?g"�.F-+�ֱ=�22H�-'-��z�[S�"�S�7�B1(R��pM��]�{���$��K!T�~e�2����FY�����o���&���b����(ŵ>��,?!=���6���.�3!TԳtʠ�!tTK��̢ȬT�q7�G�
6�$k���!���RO�N�8������.�<t��HB��T������!È�VC����dz��������������>UJ��56�t���`Eu�|c~�+�	�`�1���bBc�p. ������T���(ļ.���pʭ�a��&�z"3�wW��C�+
Ѥ���[&�4[����	�Yd�!����X�m�H7�'9�J�������~o�=�H����V#��m�8[ �&�4�!	�w�"_]��rKſ[�_P���}�����j�
����t�8�ҝ2fM)�8�et~����Hd��blbY�ӻ��_\k��o:͖�fŹ���ͪ&u�dm���e�t3��g}�
-Kh�f����4����t`?��N�n't\�� ��q=y�͖��PC��\�J�|g��k�铤�0W+Y��!!����?��������+Z�Fft���3c�S�r�&ѮѦ�-a_w�u�bn	�D���
#���%0hF8�����;�S�P�)y��U�j4��s��H���K�.b�Pu!���eH/��N�^�Q2^Tũ�-h���sp��q�Ƥ	?�}X��D�!&��i�2*��7[��\����m�E#�[�Դ��ⱷ$|)����l�gvv����T��f�8��c!��1�r�8����j�W�:����Zp#Ѧ�SS
RZ�Qk���u�V��e�W�_�X�/&�ºo����SZ�6�W#�+�F���l�dBB��Cy��O�^�=�p*=�+|�a?a8��+�-�����~VTB�-Ɨk�97�ǐ`b�"��Y*6����+�9	2�)�ޭ0^#��� ^���xӚ �F���G�6�Ğacѝ=��D����%��s�e�^��f��T�[�2lk-�_(��Y���B���[�L�T�+��h郭T����e�0Gѭ{�r}"?�����6�NB�4
��	��`v�o��A���O{��0�)�J_(�V/u�)�bTW��H����	W��qc���#L�k�;�3��P�OrnW�<e�e�y�U*����jU127@��2���&���^���[b��VԽԦ�#���N�h'QgA>l�@p�A�y�N;KX�(�p]����<�i9Kmx��E��T�k�:k!�m�s�������ð��ؔb���s��������������$�������䏷�3����g�h%�)l���n�$�4�-���2�y~9@�"�L�S1�y��#���K`��HE��5�:@�ߗ�1���$�n	�݋�&X�I�i	iC�򇹡����N%�x�19%C��Jp���Ї��~	�V��*ȗ|�d-���O��>��P毇pr���%�ٜ&� 0�~6=���"~��ʔ���: �0+���Uh��.���_&	��Iw��Y�+�˚ks���]]h��VX!R3;d+?���m�uq����/�0}�;�
�-��jڈ���LyA�_i[�\6�L�xs�B(�������(QF
SM�}�?���T�_�F2�[�N�J<=�n�-���K���k&��?���������l�C�"�o.B���o��I}oJ�݉���8֪����v��X�,����ڭ?6��$�5?��Gn����z�V�,^Fm7�� 6�4��Mץ��u�E�]cK�B��c���� ½%ѯ4�L�ő����T���K�a'W�yN���$-��Uj�6H�o'�ot�������v�#��Q����V|���3o��ʀyv�|$����1�
��ؔG�G��"�#x��!�J����}JӜ��R��!%:��sT4xhZ��IVv�E�;�Jʒ2;�{��%����>r!��e�OP=�X�.�ᴌr�SyaW�/?y��ȏyw��SL)[H�Ќ��c�S{�S�����&]z5K˄P��}Z�Xt2=�p����p�7z��g �em�Sd ��N���S���6��#Tv�|J����U	��'C��J�%?-$ݎ"�+%mc�a$�­T[p;�3O�̰�֥�f-��=((��=�ݸQ�#k��+�(G�̟�:֮��]T+4�B{a}��5��9�=��y]"X�s}�Y���J�z���(����M�H����Sj�&�FA�_p�J������OH�f`M�i�)���8RΘ��g�?f�3��&���K�}5{N˔,W _*�����_�=����&p/�ЉXh	�b�r51�37�T��Ǟ-������c0R��;`Չ� p���mBf��Y�֮%05,�ۑu�$�G��OZ��Qr�eq����H� B�Ӳ�Z�9x~�e��"H¬�2ӳL@��3�z]�Jd|��Z5	��>Р�������t�!�چ��>��R���W*�wc�2��q�����N��i�F�o�E��Òs�}���I��wX��K#C\�j���~+G��L���M;��F�g�j�uZx,�e������:�E`�-�)K':@Z�R6�����j�G��)���o%������0%�,�߀��>�.`"��z�Z�A�M.�����bc�kj�Vu�5^�B�F�cNFJ(n���=M���q���zM.Ve|8��d����:������áo�9�l��4	�j�����i1�C�"�$�^zlZ�������YP>�F�TC��$Z6�]{�`�g��CtS���a�����SQ�'E�hl#A����E!""�w��GQ.��tH1�0�;��r��!pZ]I&��:@M~lUR<�gTH`�}�U�[�C�p!Bw��dirQ�ʯq�E81"߄K],�T����+��x�����s ꨺��+�C����<��Y��/�m52��W��Q*����p�L�����ʘ�>deR���ˈ:��k��E���i�����i��hg�U�<jC������R� 8-&7"mS_s�܇�X�R����o�q��'3��#"g[�R����Z/�e��\"���/�K��ʗPʓ6�K�b�تyڢ�TB�V����Y�zXL!|��j��n�oEz�1Xɮ�Y?�nhSf
Te��7��\*�UP���$���w�=�h��dO�� ߕ�ɇ��_�r��#З�����|�6�k=Y#�u�7�^hH�	A��|3b��B�F�Z`�0�o A�?��{�����5��^ЎWsc��I��))��F �u�mTaW�{,3��H�N�Eb��X*�s'G��Y�0!����mp{f�R���{y�X�C�_���	�2j5���e�[�:k�K��y���U|�T��� 7�Ѣ'z�YԎ�t,:U���3�:ak�=�\_=���9��Oq�����hQR�;�I�,A!ɏ]�q�����5��� �=��/���-ȵ�Do�ZXR#Z��=�噵�nM0H(�o��������?�<_��_*�����;] �K7����'9,�}��?oº�i�*�}��tOHx��y�At7���҆�AH�H�K�vE�!�
I�(է�l��q��ĒS��k���)@����T8[Ve��E�]���ʺM<(zN<�����=�,��Nr�	ʮ��t�ԑ���7A��:q���Yp~hnC<��VH���~K��*&Ct��nlt�[��\@͆����$��,u����M�ʫ��T9��K��izث\��q������F+	�?��|�ܵ�ԗj��8��H �c�M��w�'hǕp�"as]��z�CS�Vb��XA��==7�� �37�8�A��#"��v$�@����F�}��M�ͣ!��v�c�6jS�������N��������
0�A���t�f| ��V9��������
]����{���m�1p*�.� �:��P+҅�S�r�W�N4��J�m�������~���>����*ű/�FJU�f�DJ5x�9��
����&o��y���OB6oQ��F�0,���֌��*����LE���]S}a�Ԍ%�a7yR���Mu����89H��Ī1����I_�r�&6;%m������[�W��Y���C�+N�;X�4i�����9��x�������}xpkU2yrX<$"?�`��HE���=��Ϛ1�+%����3>W ���Dĝ�dh��`ob�*1,cWἓ������X�l5��>�g����2TV̄e����T-�g��~�Q�2���z���I ���4�i�
>�O&'>_&U�"���o��D��# S+l{ӻcr�D�O�Q��@�u^ƾUO��U��O3;�1?VD�޴�P��G_�v{'[_5nB��fS�����X�I�<e�@���/7R>D� ~������>�@|��}^�CS�H~־hKF��h�,���lڃE?f-�]�:�J���)6��`�E�DF��4ރ���*'�^NCa) ��o�xvk@#�]j,�VX��8��e���sfff/�^ �r`
�F�NJD'l�6L~���J�f��_��)������x@ d�;Ω�	U�=�C�ھ��Ug+[��@p�K�H!��8�M�lTS�����͒j��c�S��Jk��jp@}�*�l�H�	i»i�8�j�<W����)|���W��9zf�����vڸ�B��4N:�ψ�ρU�д��[y0���G��'iAC�JN�\I;c�[b�ߚ 
u�_A{/}�r�uƋ靳�����v���9���hz�Tn���r�.(K�F��x����{u��:�{ �>�[_�{ ���	 �|��[[�׎T��5_���;����@�2��Uї�%�}��D�"��q���YH[;����U-���`cm��޲'�أR���&��#�Q��*�O1�~���sGE�k��S�{Z+��h��f��6�������)�,�jn������U 
Q��!�"~�u�A/��G��ɽ��j��|��	�y�IgWT@�@��<��I����R���x:��X�U�
�mJ\ӼmV�9�I�n�~���d#R� ���lE���1�L�)7�������&��/���\�7�8!�;���r�
���0�ڇ�4O?�]U����J3��IO�8�<.2�sTv}E�3�e��:�F�v��ڭiP�f`m���TW�k=��z����/G��G8 6��q�#�z���~�Ur�奄�݊�T��"�V���{*�qH�AW���n{Jsa`�FR�	�ؠ�J4��3ȣzv��eMz%��}�CV
����qX]�a]�t~6h�#Q�Pc,�I��/Pw�/
E�_*��Ζq����,��x�QL��n?��.%Q@Y��)��d�u�u��D�yT|ݹT�z!c���V3��ˠP���0&a	�?�$9t���:U7gYeU[ڂ���{7<�mdOZ ި�~\���v!���G�����d�Z.�o
䈧ꗢ"����D�盫�$�{*prُ[��=�d��)�x�,9�9�^B��/�x	U�)$�� �z�r2�������R`9�}��kx�yt�a��lgg����G-�\�#��-S�o\c�����O\ ������p�A��֠�|*�����N��C�t9��~���&�Ӿ����`P���e��Hp�6##�D^1Ѳ�[u�[�kB�%�Y��I��FY�S�a����iQ������B�v�C��O�@hV�]3�N�9C���e���Y�2U�C�7Ș[8zڲ`߅��$0��a*|!��"|f6=��#�ا�8ґ����*��"��$�G���6>)��+�E/���Qو�U�h6RY�����zLa˱��O��-�/�\$+���%��k���+�[��=���[�N:�{������Q��]u��)$/$-�w&b�z�b�n5�#�� 5u�3��4G��^� �2H��-��D2� �d4g�?���`s��o���^�F��o*Akdk�݊#����8��i÷-'.�;>c)[���B�f�ed�kz3��fso�͟BgY!��嗾�G�X^AH���4u�xsO��Rj�lD(���}�랎J��1�]M�K_��w��.��$)PubCc7����cK�k�Ќ�Z����,�u"a] �3�~_�=��I�P�lgh���o/��~v��'R2Vjjr	~m��,S�"T�,9N���c��Ճ/J^�-�������h�9�u�2)
��c9%2���F@�*�,�t߻;�Z���@�\���~�m�5�m�{Y��/�Ɍ�{�>���� 9_���V��%=���ʣ .����,\o�x��d���p2Q�+6�
P�$�>k��&�D2|aȯ�.߯ύ���r���b>��B�s(N��	"O;�t_$�c�7R5Tc�;��k��:��]*����΋�����U� h�����qY$d�ZRl^��4����dJ���i{|�H�s��o�8���ˋ��J�z_<1��Uj�SC��	�ʀ��d�N�E�U7��Ec�r��^eT�>��\���	W!h����O
�L1�}�A�8�R���fJ�7�����E�4�s����R�֔�������SfKF�����P�������&��r�c�:{?@%7~���2"H�M�F#��+�9�ʹ1�8h���2�{4~Wr�y>��`4L�b�3}Ծ�0����xm,�3"�� H5�OO%u9���?��{�7s1��n �2�K��k�{W��#-�������d�p�Q/���U����"Ԁ���,�D��!Vo�v��.7~_�V"7 �#�o���X1.1�D0�]R}W�i�Z}� � �b#bT�^��v0E�A:'��Y�*����'~����`0/<C�ĉHfe��v�O2���>�/ߩ�ɇ�O��)�QJ�5�>AO��[�3�
���PtQn������J�kW���BR�W\��X#�&~Q�)��iHt���ᐝ 8.(�Hٱ?�;�u��'�c�<N�^2���mp��Tǖc�0`]�BE6���.��Z�0�4?�<�㬵�p�6J|����y�.L�
[��e	2:Զ��~�J�>z�0䁅e�8*ϻ���>myc��D� ׆�n������r��<b]���� �U����Y4��d��c���1�߳��Y<X@�sˢqd,��S'3VzVbS"(ȃ;G�,?P%����G���P��\���E��Q�� I��.^V1���l�O�s�<2t��ÌbӏL���H�*���It���^&�vk�Yb��=���7�1�qy�f~}�&i��V�I;���j|o�$�"kvj ����߶+*���ڠ!9߰��سy�A�����7s�;�J�Xjp�$����~J�E� ����=�-ZR�슶��-ߑX PϬ�*f���,�:~�����4βcPe�9Y+���F1�Y �ր�HrMa$�o/־`}��^��]�_S����v.rT�arT���^�@1��[�ȹ�߁i ���K�c%[�iC�rC�	7����7 A��\��^����~ي[1o���:\]�T�i�S)'{\��cE2�n);C��u�Ũ/
�f8�W�n1�f�j���W�u�� �1�P���������C�gE���h�����2��4Q|<����ѥ�y�U#A��:�??R#Z7�M�e��$��b\��x���.���~�y:��u[�'׻�l�q��M��MjQ*%\�:�J���ā9\,���?�PܺY}�z������/�M�'�V�V_V����x��HMP�pS6bS�-x��\w�16}t�t���Cx�ֿģ|��m�gU˔�2/�Gq�r(~��F��N�L ���&�6�5���N��k�8�ztP�끏��xi��=b����������i��$�ç_��o6�l��e��"{`��gI�l�]���Dg������ٝW��Y+�m�BN�PA�:;,B�-���ș�8��2�@��f�e��l�XR��=b�Y�#_j�(��z��W�X��N��t�Ӹ�γv�>,�s�Bbe�t�'1=���w�2}�3H�;����/�&lT�U8E/�=xV���Q߉�
���IӚF6���@DJW E� ���4�-���G�;��ޫ�F��c3_�u�T����/������)E�
�M�3Lu�}�ɯ�A�`�sШ�+n`K-P�Mha^oN��aZ"�0�@N+�C���t�Z��YydT�h�yI��Jjݍ,:���[�P'n/pğ�<�̬�.P]���'u-���+0���5�$�Π;��۬}m�(�T�������� �e��b�	n<��P���E����_$^�iq����(/�"P�f��:�;]�����U(U����k�����۴�d��$?:��y)�
V`:�K��&ac�s�4���G߉P�f����3pE֒x�>�R�=��٠Z��6*sz��rX7'�3�����p�c*�Ǝj	ٹ��O���������u'%�U��e,�`(��A\D�'+���fY�:�he�UgПU�w6�x>������������
x�x]!i������ �U1�Hd��ט��Q�i@��GS�)�ɽz<��lj��/�'��kB[j�E2lͺ%����b&�lx�?�.�]T���Y�*����,8&�*Dp� �\J�@����IkǴ����n����d�6�Z�{U"NX5���t��@{����4�Og	�F�j]�]����`�
�^6�������]�W<����w��ZR5���l�F���/0"�Y6.��w�O/U(i���y|N����BP9%�L\}�Z2���İ�q��p��WuGA��	�Я˿�� ��o�[��Z4�[����d���B��{^�z��C��c�$�����r.�!kޚ����C�����o���T� {�%�֜ )Y��6]����(�y�q|��a12Q��·�D =����K��U�y�Š;��/���%�Bg�LwUP����Bq�%0,��74������g�+��(���KčG
G�"Y��O\z� ���������xS�L&�a�Y��oCx ��R8ۓ��ݎ�p�����d F�u�d:���yH�w�\U��*?�JѧH�J~���tť�.��Ӂ�>餧��P���\�,nXP�,��)�J%��P�N�I:S����[���v�e�m��o#�A�I�AM�x\K�R���s(��sO�`|F�����]s���#܌�(U1�s�Ba���?։vX�<0�n��N +��?Q��b��'�0�ə���j��|��r��9f���C]jѢ330sr%d�
��uǧ�և�-�x�.Ee��gn���H��K�NI�������]&E<Uy.�
}�(� q�����]��f|1�gŇ2���*c���ܱs6)y������(�T�(�%'�u�N�m�m�	�"�&DWyT�ѕ�WwL17j�"6m��܃
_���!���� ���*jΨ�Z(2NS���g�Z�ڐdA��	#f
�P���t�by��d���~�E\Ƽ�O���Io��m�:H"\a�cL�nX�*L)vr?��@��Y
l�����hn�7*�+J���cNL�Aaþ8���?�;�1̖�4�h��o��14�O�w��/?�e�7C~2�����l��O �0��r('�^��Є�*��Z��f�P�-6Y'vv? H���(��������<N�j]p5p��'�9�'�|�D�;v��(F��˫����П� @�TPH�n��4'�lK�gۥ���%cfl��@7�Đ����]�lB�<��LA�T��?,��c{F���Q��<�C���"�4���+�/���#�T�a5��B#f��?�- ��c�j<9�N��>q�`Hy�
����C���ɧW�P���p�a���I_��q��Y�Ϫ��N-���q�R��XO'����J�I��jG���!K�f�UAj�߆��֗3{�N�9�X��>0�ΐf�~4�U�6z\)���yM�|w��z=�#�R�/��K'�}`s���*�)�n�s��p/jy@�6���#�o�lU2�\�A�Q��Ӿe;�t$�}���BB�������qoxK�� P0��^�0�7Lݚ�")�~�Dy�����#$ZXJ1���\�Y�%����wǄ���E�V��]�����R��T��R^�{9�AM�4��m�}���NU���o��F	��HdcLT�Y,������#U@���m1�Bʭ�]�ƶ+Km���s���Q��<ZV��v��E�aH�)�ߦ�k���y�R���������vb���kA(s��M+�M��+�?iu��۟�)�ƲX�O|�@r�q�q���9�-��g)�AD�&�
����i�\��A\q)���&`MR�8\�|_\ՠ5��+6s�&�J:�&���W�Vfsq����o"�;I�b���ۙ������l��R�F�3�A�4#��8�71��r�"�Q��G��Do�Yz�a��y1{=��o�3M�ܙ�b�Ѫ����UW������
q,���S�v��MCd�X�2s?c�A�F`x�y=���7�!�KN�L��r$S�P�o@$�( �!ĿMJ+����`� ��_��[����c�&b���KaX^*�Oբ_U�]�D�X);^�m�?Y��� D8Y��N�ԕ����i|��E�A��9%S7 ���'ȇ �ރ~V���&��q���4��WMX.'�b������k�j���dW��*r$(�H���@|�:� )^�2i]Y  ��_]�mD�e�BC+U��u�����0�ڱ�k�2�Î���(���?*$�;���[���kKb���u)*��r��)a@(N:"���צȣw����d$}�K�'�����ŋL�^�$��4&ո�i�T'���E�HBTq��X�ɖ�6g//z��z�uZ���)xٮ�Mz@ت��,�ɂ�]�f!�^ON���Q�&�7{.YM���e���iw��6��o.t��tz*��7�D��h֥!���ɝ��
�XSxDC��2
	����R�͉�Z� W�����fzMd>Dx�Σd���y��
�Bb sKTZ�Ka�(o��Z�PX�.���yk/����+�͉, B�ڽ�!�.���4�O���6Q����,�X6%�(%Z�����Sk{��W�rd@��O��)��v��23m���xs�cנ����b��H����b�GR`#(}����x�GJ.�(c�Fq���h��إ�s������ns�ߚA�M��~�{�	��	��S%�Ϲ�KK<A����t�@�w�s3�|�?{'��k�8�3V��<ZLt!1�[i4Id(}��J�x��[�	�ւ��q�=b����WK6]��*U����>���C��0��1|�Ǿ��2,
i�w��q~�6�������6g�qBi�fK^kE({y�W��6n��� �m�_���	�EGH��8�����V�@\r�C/�DA�b]1H3��|���w�	��o�$l�:��}�,>�UH&��Wg���5('��|I֗>�9�g19/sz��~�5���D)��@q5��� �5�E����ss}D-ƶ�a�\8�
��n�.[r�峐Fg�)I��m�Hn� >��u
pt�dO3d���}��tt5����e�I[��gں1ҩ�.8�#�M3��T2:]Kv�2`m�,��-ޙd}h��$��x#g~C���?�l*M l@�Nh��*��n&z%!���;��ᵹU�����t=�N�hH�J�7Kt�?a�U�H��|�Vq�c�j�zr��T����ZJO�J?��FCQBc�8������o`�����mtB��ʸ�7��^��:9xy�ޕBA���(�<�Y��f��l�,�4�<�U&� d����Z�O'��Yx?�[�}�g��m�]�ٮ��g8k�^;�/t���1���i0��~ĪXΜvI�m���S��˅{E�5��Ag!�O�|y�
q[�2�b��֖����� ��~�~z�T�f�c���C,0�|�g��gap��V\�?��>G�h�j�*��2��������&x$-�H(l��;�gU��Q=����֖m��_�ٗlc���yZ']��pHS՛q�W)�F�v���ج[j��\�l��� ��g�awA]m�l�آǗ����v3�V=_��s6�j��<�w� ��m�s���-�a�[׼�_
�ə�H�0��XwX�KpK��{2sh�R�{���<+��
�T�,֫�R�n;?��y�f�yI5ak��s�
k�b��D#4�d&��ײ������t�t�y,���/����%X�o÷��x����~�1P˼ےk�K��4��+�
�D>P��
��2Y�G�������@��V����N#i��^}���B�u��ƶ~�:[s;١�';q�"�?��
+ҭ�=�9N5�ĭ?sO>L6BTz*���rj��F�K�Oq]�4!Vc	�d��R:գ�����tv���?B-Kc�a&l��Xǣ�� [�TY��r���][� ������� {gOA9���*��~hOҎf�k� �EW|:+T2x�܌=��f��A@��n�'A�4h�ײ���栝��V69����^�)Y�[Ɣ���1����NSd��A��i���uB�����.~���lb���~�B�P7��  ^'�E��wdIF<Gb!�����U�)F����W'�q�H���5O�#�Xݢ֎����hl�P�'d�ŏ-�竰.h�v�~���A�=i�n���]�Bd��|!�3\?�5�1��(ft���:n̫�.n3�ƲôĲ���я�"�ˏV��H���r��k@3�+�g2AP�K<'An��]?�P[���;`�#Ď�<�S�>�`��(+��R���q�8�$q.�bВ@���,0�g9�"cx+�w�YFP�_�a	}<y4UT����Ѧ[�	P�2�d^�,^�C���j}?/�p:2����j��nt?��8X�5�-<w�IqNd
R�>n����zR	v]� ^��Z���c��xT
:C^䂳�rG�R����A�,ޙ�d�b�J�[�O��d�$x ҕ�	NH�Iϛl��DS'LE\���s켝!�S"��<�d�|$�a�W0h{V{��5K���<j�����O>%�%^�6
��+bgx��}��:0@������5����+ķ�j�s�ٲ�~~G0��<��D�SqDђ*�g��U�h�m���O�>�ȻXJ�7mJP17��8��`,�ɥ���64�O�7Z� JQm�5#!��5���f�lJNp/(�r Y�	�h1%Xiv/_T\�M��@7�C\�)����Α1X��W�絬&��0Pfy��IY�?���j���4x�ynߙ�ECzl�=����`U�?�\b����@�nO�>+^�@�/����B	�zHm,���h���:�^�VZ�����Pg\mҍ��@��8m�B"g��I��O�a����ԓ�/J9,�$�j��-���ѩ+����I�_3�	+|�n"}i���4|�̠���Py�L�rٓN���i���3��q����-<�./�Sra{��Y��XY>l�G�m�p�7��-�l�f��`'�\1���Z�c�:��҃��:Q8�y���Sj1��}E����3���￣��J����4�0%k�C~�Q�g;Ei9�,�����-�K�[A��{��B|d�ɺLēf_�,�Z#���!BEG���Oʾ$p����y�
g�`�x�3�wz�<�[`��JV����8Z�����.Hn�;P��?PFѢ��%�>@��ZG4p,�� �&���jl;6�1J�o>:=j[��cF��6�c�F��֜:����9���bw
���@q��O��$��&{w3@
�L7Yt��F{/o�
8��zQ̦�0���1�P�(i���R���y}4Ɔ)��:C�\�ِ������̗7��vy<|u_��E\�n���1Iל�6NBu�J�r�yw�Q?'�ӊ���g5��
�
-'&��h_1�*R���z'f�4v.�ts7�F��E@���i��l7y�CO2Wvo���vZ������L	���*O�U��_���8������++aC�<Cƍ �*^~��^��C�e�C���l�E���ۮ?� ��㜛��7@WE6��~�O	t8�0.NV��̪n�������j�f.y�W�߾&�m=D#�a�@é֒�36���O�"J�I9$��־�d8Ո�g	 ��5�v������,�E��(�l��APڪ�K�%�w1�"�ۥ�[;�0�[7�z`F�˫0m�cĲ����Wn��Bz�td�$�2���n`���-˼��6��9(���^;oE�=�#"�ȶ��ܾU�96����o���N� �6b�ʯ��!��b�e���� Ar��u^�#��L���d�21x�D�:?lg��6PCy����ẑ.�Uv��
|g��-���GMEL^�l�G�D9�'�M�}�0XN�8����G�R��I���m�,��}~�C�m�w���	s�U��D��#j������;���2_��Ҽ�PlD�b7�0�$�Μv�48�vP�(<����{A�\D:U}I&wK�[�s�S�C�F�§ K���B��+[d��+lf*��r<l��.q���}f�Jz����6
~������'�v��7Jد�x樫?!��Uu?Fe�6+:Q|#T�q���?�s�8U���q�֚�_'/F�>FY�l�r���1�6efo�sa,a\��oo���x�����w�a)�'�?�xKR���|����kD� �+$���^w�M�g(��V����b��U������_TNb�h�r��?Ҥ��X7��j��ß|7Xp�>&	��fF�+��o����'���K��j[��q��������O��zp���܈��f���-5�΂���w'r&ۺ坑�Z)cm�giDzq�u�<,�_W�k�
��J���Z���������JX!'�6�Q��B��ߥ�D�@�c�����a�⓿���*f@
[v/d}��fMbq�j������	�f)Px�k�X4��ڷx:]N-�_�ے�>��ng�QH!��~��B�=`e�`���8b��މp�g�sC�pM[�8�n ���Gi��=C�b�'�����h�r2w����5��=��^݃D�P
�dm�߉D�a�k
��l���ZD�u���J�u8Ya���0�g��j��8w;�5�A��������Sc{�T�"�\�����-�Ew.r���`�I 7,���aa�<(���rc#��J=��a�B��C��ƈ�v�K��	p����k����/��5�A}Y��G$��uKO�Wݼ����,�ܱ���c�#Y�F�n(\�c-�[CB!A�-��b��G`LkT��aW'
#+83���U�X���zH��ʄ�R�Q҂$s�H�V���hs��tv�Ɛ��J�Nu%������hP!�^����z��;g{��30<vm2(ni���<�MY�x�<]�ԲO{�z���|6�Op�A�{�±��᳖/T��*ś�eM*����fT�JU����@��q������}����y����R��mI(�v"Z'Ι�Jz`����]=m"���&������W���چ�8��2M���u����{��
@�{h/�rӤM����ֹ�'Č��o��DS]��?	MMu�j�w[����к�`��V��~&����d6������t�{�ĩ9@��m�����k.!��u!��D�Cf��F���\�e3�)4"�J*�Z7�yʎU�c�!&�D��a�x��C	��韨�XՆ���{�����?}���?6p+$p_�ճf~R�E�3����0l$L�MX	��\��5��\��L��UNt��_h��(`5�&h�1M/�����q9S{��g������J����p0kP�>����'����u]�o�����:��
	�L8 ������j�ڀUXJdV�E�[�}#��P~��ȷ%�/mȕ]�p$��Q	��O��ve�vp�Qin;)��z�����T�Z(��ۉ������s�_���X�O�+�'�Dٛ&��\���66՘Nۄ�Ѕl�rwR ����*IB�m_l8�U��Z,��g�����/<;��w�IV�k����~�9��ݽ�"|M��"!+o���CKq�Ic�5�{�>T�:��aY��%Q�Թ��Zb�8�!{�	����\�}�o�jc���2=���p�|H�8:���O�o�П;*E��N֘u8��Ye��r`J�Q;?�) Y�6���'��~cZ��i�}�2cCK�P�ݔ�&!������a��IaR;OZ�PǙ�Jw���xEı��U�Àu���ԘZ��≫��(2m������S���o���D��T�d�-t�H���Ud����zj�~H���Q~�9"{���E+�d_H������T�|:�k���A����&S6ap^�$��PV2	�]%-�$P=ۓ��H��O�k=X̛@�����i6��'�Z�/��ɗ���違�(J���A���W|}����j�(��A홺e���~o�|����zWL�+c5�?΋�{� �З�B�ċ1	q���^͍���S=P}���������7A"���)��%����''n��h�R�.���������x����u|�DS*��}]Q9�dWn�Y7�R"9��=����	�*�%�^�_L�EA0j��)e��z�[��_��*���M�l��j%	��1}�.W���Gu��rHV���Y8�*�������d��EMppW\�qɻ,za6��5��.�y����}�3�9�W�;�g��)�x]��`�����hV���D�h&����� ������u*U �*�k�P�V�䖅���nX�������Q���+�\��+P}v�(�2LB�	z�6zj97'�K�L�˄���V�`�\�쳫ˤ�¸�G�@:UGF����'�hvUڵ�n<>^�7�"���޹���	�$!>�P��d01_�q!Iϲ+�Ġ��gְ�@��4J�L�x�8}��r�SBLc_�8��F��h�B�]�5a�
�
v�n����Q��q5ۻ���I�c7;MW���U����Ml!�!۝Sy�7�I�])�kP4���E�q��y��*e�\Ί��T��l��y�O��ڷ#�pIQ�۪{�z�q����޲3Z��������@:�9�Y�G�|N�փ��	�A$�f.�K�E@�ev����F��=�~bs��vӉc�u`��Y9/v騾h/@�ZT.���Y2�p�	o��8�+k��r�#U������>���'����v��J�vu{w+�D��j�� l*7�<�.�\�pi�mC@�b4�ۖ�^-+�y��r�+���@���<�i$��W�V��;9oL;����CDq{�C2��oR�cQ�g4
�l�W�b;��P���q���.��NŘ���,m7tNa�WO����sw�ۍE�z�l��<{^3���8 �+�g><��s��~؈;Be9tn���������L�,��b ���6cS2���|��T��ZKFf�((�g*C�i�+�Xt7�~sM��
�v@)���>Dm.|6m7\�H{9�����!�>�kBh.*w��F�~m���m�ͮ�US߆5��	4��F[�߁�F��4�|vC�*�r)��=�rrcO��HzhN@(�)�[�{�%�˲��b�Oq�#QF�L)[�� �Qg��C)� 2�1,$���&�c-��|tŜ1���g������X�RPH�����?�RF6�D�Vf?��F�I���wg��ſpM�ב@���>��L�x��g��������7߄����%~7锃�=�	�%���Y2��������I[�B���/��ɪI��g�{Y�� S?vk�pv��ib����+�v��D�vV�;e���� �.����l��W�sӔ�T���8L��ruE1 ��YE.Jp�T.�W3 ���_> 4��ΫK�z�̢`��H��C��x��P��I�۫[������x]e�#��w�~DO�qe-��(k0�B�4�5@S?�Y9��}C��e�hx*�ȴ���yN�A7Vs���N���09�o��{�U$!`_��~*�q	�|is�F����P�ƅ�r�
2	�$�m��'��I�*�e�'~���	p�?IH�D�����d���RF� gů���H��h�1��$
9�X�����U�����
���Y��\���� /()�)=~yL�}˹�H�r�}��Ȱ�YM�����/��Z�޲�t�G�qxb�&��=:Z�����J��22��RI�j��G@�oeUSr���!���D�Q=|4E;�tB��g 뷝���Y�ΓS���4�����6�,|�hn�v2H�W/m_�-�&���^Dz\���e	�p��^�� 2��s#@c��2������\�+X܁�+/Y���4����0$^eq�.�tN#�	�$Vb�vҀl�+/G ��e���ʶ�G�?y��b�F�5�9�
���sO����o�S�F�*D����6�U9ӑH���r_jH��Ay��?��rR�_�>~ݚ�>�Q���C���;�8�8���U"��o��EJ��.�3E�¬��������`����y�dBx�e�4���R����dk���ZGx�0ID��M>e�z�t|����P~��<貿)��+ڲhj��ҿ�5;��W�g���=q�0�� ,��ڦ1��+@#a�g�M��)1^�	Щv��:����������.6�y�X'����+h>�{��e�E0�+[xK�mP�����G�6�3����W�o����Y��7�u� ���Y�u�@L�m�u�h�m����$�֮&��ޭ�k���w�/`Ǘ�D"U�����W����aE9��D�HF�Ǎ|=)l=�̺�{�y_h1c���z�bp1�wO��&6M��2�Ogvpn��,7��XNRµ)����#��2�
�L#Wvg�So'�i:�*A��{l>��m�@������`�	�.���Z纁1<�b 6�pY��X�icE��&jqk�����&��ϟ�#ɔ��*�;�������k'^:�"L���~j�d|O2��a[v����S�C���y����O�Z4>�N�{qa�2�3�����qMl`���y�x�q�ْ��m��o����eq`X�#��D�1A{������+_��K�����,�gi�����Q2L�Ct��s1��\ͬ�>M:�kn�c��)�w��:`�ǳ�R��>�G툛l�`��sZ��"�yTh��\d�y���J��nUb]\O �X��8��T��Ѻ俨�4b�7��d7
}�J�꽵ZEX���,Os|��W/>1ߜ�a�aкux7g����Gx��2�<ᴢ��Qx��±��|�SIl�� ��tڊ{"� ~}-v-����w��_�fh���.?A�Zn��)n����0�}Fa�ߔ�:	=骐Mt��*�G���=���5[Dr�jX�nu�ᵙ�h
ms�i�y���PD�� ;$\��=��[q���O}���x�����!�� p?���H5�8P[M��6�Y�U�3F�n��}��od6��C>!���":7����Ni<C�$� ��B(�d=bmA1��վ�u�,]2wMX����
�
D+W'��vi�W~�-v�B]�G\ц
�mV��e�2��:�	S*X�?}���-4�QK�ybM�v�讱��W[�53,���XB���/dI2�е��Z�G2χ%m��FYa�����	+<���s����s
��ޯ�˄� ��H�U;?�4@��7B�?l��&���՛�~���12v#i�z�@<�[�C��N_��d���[�B����y
���#�����ߤDz�T�_�0��Xyr����ؘ�B��H�8�S򧺚���Rߴ�I<l��5f,_����s�"��:&ۜ��2����HHZ����9��|*U�&���7�z��ަ4��K���W��%hQ7w/�#��m�4!�u袇N��̍f��
x��b��ج-�����M	g@	�ZOi��-[V�>�4ʟV²;,u�q������d�uO�j#n�#��)F��Æ�J:�y�ȂOX�cP���{�1|�j;gհ3��q۰j:I�j)r�t��Af:�s``���i|�؜KVF�^��g&hU5v�b�za��߅�q�Lm���s`
�2di��[�siX\�����|篚���uo0�p���cJQ)l֨r~��'Kݪ��J�������'<�+�bo�Pفw�qOah��R�Sg�@�c[q�U]'*�<�z����A�r ����T��1*b�?��v�ڔ�W�
1 N�:\�ӹ�Z/)� ��K�ãБ�5�H�j~�i/E**&, �t�B�#��)�H���z𽘰�K�/�m`Z��n�l$m.�����05t !���(�)v���*x�
*b{َ8� �C���B?��iT�{yǣI�Iբ�M�x���Ĉ�S\����﵎��
�K���p�����{��Ub��%vH�K'��I�(�Y\��N�]}��E���,�ѵ�f�?+`����r&{�VV�A"t���*�s�!���P��^�v$�|Bv�4^>��X��īwQ�=}pQ����3�K�[��A��{ү��c���3nެ��TlFJ�ȥn�{n��zp�#�	F6�����9E:!�-�ϯ�fXWL�0�7bv����Q���� ���̿
�e+;(z�ܫ@��/�>"�/��­������T��]R�Y��$�.�r���-Q-" }9���9���KӜ�����A2�s������f�z��mh���sw�F1%L�dF�N\y�y@�R}$!߲�b�]��$�H�8�8��ߕ�=��5%���t�;�h�����YA���'��)Q�$qO�[��� ����&;9>3��0KC���C�����~kS�?-�P�%9"�ݯ�:�"�X�X7��\��B���ՐEF߱-���n����{g�+h�`����_�Ev�m7+�(���O4VV׾ow^3����o0N���奦�!��.�]/���~m[h���#��z�nH�G���h׈�N&��:*Ȟ|)D\D}b�A���.4� kJ����W<�v·�n�;d�d�$lT�=�.F�5�H����A��$R�ګhf8���x�E�a�,���k� ��77�R�ٵ�,.�OD��)�иT���:?���c���a�,&с79_�����������|��W�3,T�����Om%%�n �J�zϷY�'Z�9Di�9�z�W�ڬ��dr��͓B�IA�c�=�u�CAh��N~��1|��^5�(�"� Z��Sa*��N�3Ӂ�V!�'����a�_l�	��Zh��s\��~v�� &�/ļJ��3��F��&n18Zy��W�t-�j]M`�Hs���%�s2�h���d�)ދ�0��|<���ք:#���νj@���u��z2�&pW�OǇU�S�9���5��q!v�"�S3�(1g���c��y2�Nހ�L�!����}������OJX�e�w������%D:��_���p"�KI�^,���EF��eg�'���4S����0�y �Y��ͬ���yF��f�*'b	�`��&��QLSlk6_��=|�_Ѣ�ԋ��O����E��)�h��Z�3į�Yu��v��H"�w=���|�"n��g�?�XR}VW�}>���86�M�l�y��A&��:�ؿY��v���~��{�&��8��%��9��L,Ee�~���7t00���3^�y{�7͏8�v��[E���xxD�:P"�3�BvA�:y�P����I=s$�l%��|��p�a�6�>�P	6`�*u-�O�&�Z(�'�c���mO���5-��m۠�pNlf��vB)�N6�xv�\�N�η��$�j7:�CnnU�O��nl�{k�r�B��Oק��[F�-R��A����f,¼����4�W�j�����c��l��[x�H�K[���!%hΛ��sͻN��N0��GQr A&�FS
��х��<V_�����x��i&������������4'�cF�`�5�Q����.^B�Jr��F�v&���۪��҃�>�n8"�`|�4ݧ*^��7)0��b�VO.�Ǔ�3�"��P���eM�jc
��QO�9��A~|���*��ۣ(uP��&ޅ�4sd�� >?�(�$Da�.��B/O���'b�o?�t�2�5�ƽif4��.����o��`��܋���T8W��Y[b�(�-=�&/�҃L�& �AjX�إR�O�R�ٯ� ��6�W�K]-��6�2�`�������-@e�X���U�%����g 
Ҵ��H�$]��2��N[�sw� ̗�Z_!N��֏|3��UK,��HIT�@�+�����������z_�
u��	�@}Y��L����*���8�ԯ�#��Ϋl��:��%��Oa��q�X=�B�5�94B�*���e����^�j�T��/�
��>	�^�t�4N�<���i�p�-�{>{]	�J�����qÏ+}Y]���|�`�H��Cn@.P���y����A%XDT�s�B�?���zm� ���w�`T���ɟSv��6���b&ibc䧄,ȔY��aT ���v�w`����>��դ�@o\I�׵p�+��!j7+�ki�����'�����H�U���?�נ8��H@)Q4�D*�������+r��p�$����m���4�ɍ��78���#|.cm��``�(�zCB%��(j).�M�TCd��>3�ač˔K�?*�2|L	�0�;fΌ��ju������|^�(*'��b��j��O�E��r�Xg���?������M)���X4��`�v-Y���%��'w�jv|�#�۹(��>J�[=,�NL]���=Z���k�c~�0>9ŵ�Ɛ}rUtXzv2�ec�k�y`V���&b��\�v{nA�	�����mv�3^�"�	I��J����I�aqޢ4�I�G�_�N���Z�f�Ѓ�����5��4G�k��hslv�F��u_������"a��9/�WQK�&r�=@	��&�{1�-0�yW�X&}����=�!b>�>�ې�����<��9:�]�_��Q�B�:f�i�}3�z���8�n���\�H�M���.]���`~
.�I��{_iێ(�|�;EkK����޼���0�G~�"�u����I��`�ʛ4i�&��N:�<r-�}F�IF�¿����_j�
���h۲-�RzNɸc����s�Ά�@�c�f�]�)��a }�~^��gʿ�H�����
$3v�@���u��]M�.F �/��(A�Q���!k�7�!\�B�&���H��^�b�0fo"�H�)�1����iޒ�bs>�Q�QY%
%�%5�m�5�����VE���|� ����Tcx|t<WZ���@WV���b*l��n�%я�_�ÌQS��)}�7��&�vo�,=sDt&.U(ҍ����
��[�53���[Xw����,�~����"kѤo��e�v7m��!�XT�w�n_�a2��#�- ��1X X��bXe��3_B�6����P��D����$��(e��y6��1);�߄{|,V��4B��z��x�L��Y�m2��`G����>c��Pc~}�]n��v���"�>���2�$���q�EE�{�Cф�'#(!���ujAԙA)�L�ƽ!�^�'���_W���ذ�1���B���
�Ѕz�&��d�`n��W��aP���'eċ}^r=GƧ�#<Q[t�4��0�EL��>�j�UH��27خX��������+^����E鲕���h��Pǭ��i��[	��RB�Sc,P�UD�k#l<���d�j?��҅�	�R�֕�`p��`7 �MV���̠ע(���\rrz��K󨉢�G��	��҂%�
���2	�P��<�+�td��uC��ZNp��޷8�y\��7c}�0��4�)�S��y�?n{�܃R互�M勯{+�WuI��3��anM\P2�-�y�Xiz�`�Bv�w˧X�a���\H~cv5)����qH���(�
0��C��,z���X��UfuP�G�Ƚ�{����6�`S���x��N�ӱ�ؐ�Z�[�τ�VL�DK�MUmC�+5C²�59� �Z��F���'�{y� i��[Җ� j�� K������D�*[|�IȚD������A,+��χdшa����/yL����7�� ��e�z�����
�Ny���Tj}�1*�ߝ���[o�kS}��iG6F��ͿQ���1�uf�	���K ��9�Lr�N�G�_�0b�K����P?�.)+�"+����i<�s�E�ޟ�aŻ��*���F��bƤ�r 3�`�Ɓ���G�%�nH��_]-��Mp�~�z�}��٨P��#�������%��/8�s$]f�`�vzA�?���1�k�*~��"��N�еON.'pF�*բP����N�%�v՛ܲ@x�O^XX�K$#�s+�7�C�ֽP�k4�e��ه9Z���U��s��U��+Q/�Dp8*������l�DH�ޝs�+eb�Q�^|�}��S�J��xm��L��!��O3���5}��"b�F&��dF�G%���o\d�}����{˼��tv5W��Ǫ	g��.}���<!_�a����D�D~�P�>��M�v���L/�F�ŗ����޵!ؐ��\	m*�(��
�����Ωi]��aJ�����	���H{���ɼ�sMWWT�%�K�l����K���ҁ��J�3�O�H��Rd�W�=���DĮt�ն\��~D���g�8L|$+x�!������7�ZU���d�R��$�+�!oh��d��x�+(`bhrR�;"����d�M���9��gȂ]qh,���(e供Gg;lI��;D��M#�<�^����P�/y*�"H^N�Oځ�p�1�EA)�&��3���ғ��U{Q�3��ʛ��x�+�,��DUVL�)�%�bX��/DJ��;���Ҭ�O��� ��kl��C�Um�cB'��Q_)?]Yq��e6Z���5e$%��f{Yy�I��M���>�\/��5�K �
�s���&�Y����f@��Z�:�6'r�@���dc�7���0Џ�S� ���*2|UtjUR^�� �/r�%���24�����i�Z��_lr=+E���m�>�3�G%��.�z�@�l:"�T<������ ��K�3�Q�it�\qЅ	��U/��/��%A�+���4CE��6�:�n_�Z7��qb N���l��e��@xNō�mJ�n�� F�IU �:_l�?�*��_��^D�O�ؐ�[��`���awb�H���MPHQY��PrZg�3b�q��Pم�9Q#�q�����cм��� *�|x���i2삆{
���4�&H;}ކ͂��/�5�IZ�^� {ܫ@����.�;�7@fO� �i򬝕^�'��m9H=,`�Ⳇk��	1/ßhp������'pU���pm�vȍvN���R�В�=��PrW܄>�G+])�&���H�+��c:
�&ۨ��zos��G2��/�̹�+W�����C���3����:_����hAFܬ!��|�YG�� ��ߊY0�!/ �SG���)��mG�LB�A|�7���D�,v���G�$H�F�7V����y���N:�S�Ŋ�'Ny���pw�&��nӁu�x�D�)(��͛B�0R���y����C�u,J[��l�PwV�O��|&�?q[�q� �p��w�ݶE%}���2*�lu\�cP��7RY�����0�yF�U��p�CtO����}Ώ������t�-p*��cc���Ǥ&�.�w���L	�'Ps��cp��%�B`h�07x�E����x��Ș#�"���ʝDZ�"�w�[�M�<Ż鱸CF��&�l�x7�"�/�'����R~i]2��sv35>'�쥬-�x:�)�)eD+���R �Em�fT���w�&%K�K0u~��et%h��V��2����"�0fa����� 'k3ڏ,�(�[�32?���zM�5b�m�Z������;��ߥ�C0�40�mn���4 �_P1�W!oW[	-Q�a(�Lp4q�S<F�p�o8���|z�E98y���&���6-=���j�>)�����8�,��a���DY��]����>F�pL�5�wkx?�v����)y�|K��f2�ߩU�H\�~�ȿ�WQ��dã�ÝX�yAV�D�p=���W�z��)$���j������^�`)�'4)�F�/�S��	�^��}�[�g��� �O<[�'Q׃��P�U��#�H;�T,�u��{\������a�ƾ��ɜv8�m���i���׼�[w��(.(�/pH�6�t���s�Ӽ�OQ`=�JQ��W��4.�'�G�=���byW?�-$��Fg]K��uŒ�s��S�	]̗�Հ)�������d[��I@�"D��;�[�9�W������W1E���m�Z2WgǭCW�SD�|�x��vm!�= �5⼧;��Z�qx������"H�t�P�g
�-�!�#�:���fd��Ù�:�7��a��JXʈ��^�t��⨂�7��׈�s҆@D�
-�xRE�O��������r�_PQ� >��{QB����#Q�����Y�Z����{m[lx�+Jӂ�7���'�k0�ec�Aow_BQǚ���"\Y`r�����tk���%�O� �43^X�� ��euꦶ��;{w�����>j��Pm�W{5[�:�ͯ�lJ�e�fO4����gq��*�u�AuR%���k��O��a��T��К�S�cXH��5�i(�[˴U��a+I�񤻴׬�j`�*f{A���M1�����dP��+-mߡ�~��l��E/�i����C����O��8��I�n? �Ua�A��)�?�@dr�r��&�׷�^{�f-Ka��vN��!��q8 ��E���H�ھX�o5�m(�, ��%�F���v�%Z��W�!�jmwa�o���6�Ċl��(=�L�ۢx���"E0���k�Xgc���B����8hEۮ�t
��6����zQ�Ke9�W+*�������Z5�gK�!fh[K`��̓?��
��O�V���V%i�O��q�t&�q�Vf�?^�y�I�kMZ�yGX��D�i�UI����*G��F�ZI�$}��kYV\(Y��A��u\8�w�HP��)x�β�%SS�b+'r~��|%6��ϯX�cL������=�j����4@��!>c��cZ^ %owY�����B�&���=�l��oi��s�������	�^17F9�F� +��K���I��,:�C�o�Iy��̐j�`J_�b�LmM�g��A!1ɐ������%�k�~\�p}��%$p�Pj�m�������'UԹ�3�vȓ�Yc����«
������� @�>�s9W8�*��w�,��a��Ȧ�뎑�VƑ�����Vv�/�*�R��s](�<DF��P:�z���Ap�	ԥs��?�MF�z���@���	�7m��4��Q]j�֎��@Ry˥'`�=1�����*�G���=ܗ�:���=+Ŝg�J���%�hmH}�ej�c��vȥn���zs%`�m�P?�l0�V�fںg-_F����Xp�!H,�\��N٤��;�|��u6'��C8���ܘ��G�/���g��	����,]�RGg����a�=�]�%]��0nXM(��d�4�T�@�EiB�*��1jrX�l��q�V3���r:�>蜛ל�d�jC�>�8M��Kd���&��m�A���V�R��k�N<W~ھ��a0�ZV�����\��;�fY� ��5��K@���$�������*�*�X�d�
<��ǣB��<c���R_[%���;X�G�u�2A�єݰ�D��;W��䇖��@�'Oe!_5(�p�ܕ�өK�C���F)����W
p���h��K���D���5����Z�/��[5n������Mf؃XA�)�'�ڇ�@զ��źF���Mʦ�plK�ě\tn�����l��{|��_Yb�r
2���؎>�p��N��n�<�/`c��4�r��Z8�����1�������O~1��l�Ԅ.L������Gd4�%Ί�=��c�ƙD��d������*�Tb'cb^�7��I��ٿ�����NQ�$�0�Q�.��Ƒe.s���l\W|±�L��|�[%���#���.�Ҭ����{^N��3��`P��`Ө����Z)|��qآJ� si���1C���sH(U�ص�B9�a����;�h�YjA1Y|GH���h�5:M�fwΈ����H�ip���Yu1h�J����&G)�;�W�L���vϸ��T�����_SN���MV4�8o�[Cb�ݹ��X�t*��d�~hs^]��EhYs��1��3H�V�Wϐ ��� +�ִ��@04%�mV���ND�0���
�񑱞�y��Ę+�rj���;�MDX�+�c+̫�ϩI�ʃ�@��
��M�+/ww�e�|i��w�V���=�lLg�	X<�s�(�j��K��d���Q\�4a����2�;\˴uI�:Ć��ٴ��C�}m�d\߾I��jG���&����~��x4���<ʭ�ew�)��B��i��|����b?�:�/>j���e��q�8���X��zB�?Z`w�<D2$��$K�`���X��XV]h�s�ۢp��f��څ�+n{�����v �d��f��ʰ�s��Y)��l^�`k)������Ո}�Z�woU[`.M͉	VX�_ۖ��' �a	٦�ء!�\%t����[�(���ljLNRa��'�ٟ��������w���� ��VY"d��E,N�Ɉ�80L���K�e���	c�ϖ�5R4Ţ��K������g����Ș$���Do�]�4��hè��H'<�_89BOe�p�)��E�����t�M{���G������O�2��B�`�l Ѻ^C$�Y�Zu�s�(Ty�I"�nڠ���q�a�W�G�*KIE��J9��,ZΥYZ�s�#b=��~��7h�u�]JXy�T�Nq�>5ǽ	>?bń����,!Qi�"�u=8�����|�K�|��4����Iq����;��*���S_dg��5<)��)K �u�3ǁvp��A��k��yg�vT���#s65H3��(�3I���,l��b,���D�$H=1}�Ʈ)�>��D��Ύ\����<��9� c��A�PB)�	�(]�[JV��\�~�H��k�X�b��L6�ʬ20ꢑzǙ�k)�.�zs���4����n��/�E�o|Uˑ�ڝX����G��L-4�enz�
��t��'��kzx�#��C�i��O�n��i�8�?
f�D7ǒ��GGU������ޱΈ1����)+���E�c��	���҉�`��+[��)�a�	PL�>�M 1c��d����=�T�H�w�+Ύ��_qi?J)�.���>(���4R�ѡ��I��`.h_v)I��
�����qYP`S.B�l=iK�zzdg���Y� �H_U��L�G3h�]^�s����t>c�3���H���F�d�l�d_fK���Lp�,�²���ܵ� d'7��K�eWɊ�=��� �M����������S��Ly����8��r�@ՆG����N(������r��Qߞ ɦg��p성�W��;���}�,~<O�q�F_�K��B^�>ࣁ@m��2�ؚ)��?W���y=<Q��.�o���[��kϙ�l�AP�Ֆ'"Ԩ��� ����:���*��B�_��KJ���EVJY%y�w��X�[��Xt����7y���y�+Hd=`i]c�\Qˑ�P�r3S�h��߀i3�0?le��.r�zO�\8_�Ac�vS���I%W�4�vc�@�p�6�g�I�PR{T2��w��[�Ĳ�ߜħ()V����<��Y�l@��%6�Z����ݑQ޹����U�bc?��OC��H�F��s�&<z�\Ƣ3@JZHZ���B���sh�V�܇�9s���A�ͱk�߉Ͷf��H��||)������2e�F����,�o�*�Y�)�h�qV�.��<˗sզ� ���<�̗^�	�����5G(nY~���vL�83b��FХ�^d9���k���xY9�&� ]�H��wNVc��d��|lðlp����tg�ĥ-8���uO&f�( �B���E�T�@޴8��49]x�n�{��'���)<�DlC��.�']�B'�R2܎���U��6���%�J�X�!�-��7>MCd:�Ƹ����6 ��WmZķ��U��'E�I�[��ck�ۨ$�2%s��V�2�ԣ��e��i$��k�j��1ؾO/,KdB�2G��TϤJ˞����J�u���&���	-Zb����g�,oX[����K�@�nI׫�<���i��P��I�:�/E��~e�����r����uϜ(��%C?.��~�46��)(GA�B����،C*��q�L�8������O�3�F�Ƴ���N�(�!�?g�g�i�[��.�?�aFQI�&�TG�7�3�N#[̾����EP����G�_�����s���]�Y�]��ZN�m��y�݋B�06�F2�T�S!X����a�|%:�B1(/^v�g~4�t0�U���a%�7�G��� �3�O���S�VvLM*���t�,�˽�e�eG�F 	Cp4����ݮ��4h��#瀻��s� �U����a��I���I� ��'�ƿ&�W@��V��WX)�9c����Hi4�(O�)g���W�5����g��"���?���k�d� *���!Teۼ;N{6o_F*/msm#6��C��/�#)(�lH����;���Ў쵋9֞� �m#1�^�>_`ə����b����-H�C��X���x�/�L#���	�{��R�f���:̙�A��"��db�<_�O_�'�N����[:qxG�;!��ć�#L�7�>��|��_Z"?�	9��+!լo)����5�n7��/�/r9st��wQ�3�g5�q�	�Kk�����H�.���.��ƅH;��Xe��bI�~�C:����0�>B�H��U�VzЩ+���Ľ�Q.%ޛ��#����E~����/W���ę8 �D�����c+Ql�8
�D�_yԄs���ͱ���VQ���t������Q��������;$�Z�F�2���D�+ �O)g�	���,�y&C8m���ѱq$�m���~�����̑��|��<|-�큋/��8�S�>�?�OT�}ୖ_����tr��Ʃ����į�<�@aD}��7v���(��t5��ޏZ�V�f���&Z׾�"Κ�K6��nQn�������w�0�ūܠ�䤬4�~G���U\�9/1�y�W�����ա���B�b�Qcӭ̲�y^�|��+��e����/��*��	2�*o�Y�0�U�\���t���yH��mn[sY�:�&xr@&4�M���
X"2�� W v3����mI1�PV��N)V�`R�4�L�� �Eȼ��S�)���NV��G�X��ʝ]�,^0�ٓ������O�*.s�4���Qy�Y>G�xl�W�F4>��c�O���?@gja�Q�,�
�d�%׼0�W���Ib�"vZx=����H+np�a��1�%��0	�[Ӡ�权v�"�3k��X��DSHf�QrfYW�c����8�υ|V�>�>B�An܇�eT��
oY��י���ÑkBg�dr������O%���t�,D����b$S{'ڟ���!�F�	P�uJ��'6XQ�����?�A�+`�o�H]#���hX�!8�K�?�=xn��?�&�x\vpR�*�}���nn��lun(����35<5󙷓��y�6��$yu|V�mE�T��d���+;2� �w�Ro�P@4Z�7���l��2����6R�0E��v���)�f=U���A�pޢbDW��^Y&K�s6&�=}��	����7|*A��3�Q+�O����<,�(-����8\�]����E���.t�+ ��:�:�S��
+���G#c��T����`��qu�2p�i˶Ēu��dP�R�.�u|q?�,����M��~��b�!L&IT���ǌ�&�Ŝ��y??��Fc	0��ڸv��t:��Dhy���EU�܋G"�|��~iǾ�@)sL��p�8�5ղ�}�~�3�0@�ED��K�R����(7h��$>�7���A���
���kh_1�=i���&{�����7�И��m�&�~r 6kr���x�z�p��b�u�Z-oZd׵�ȳ�~��PΌP۟�=���t%����-v�J	K�cV8�_Ϟ�=[�M��(}�I�Rh�U޴�K��d��h�QdFy��w
�z$��g����_�5"}�i�9��3�i�MRL�l�~P�X��ܦ#ě,�)������3H8���Е��4G��ƿd��!,�~\�Z�H�R��c	)*Z�/;+����sd;�ص�#���� ��w��2'4S8�{�l����/h�3����ݨ���ig����?E�q��2�DJl�fHtA�0'�Z5�����I����4��"�R�UP6Pf������ڤ�N(�K� ���!:잖#�2`¶�R�`<�5��va5b5�1��F����p�T֠���S+Oh`ފ�P�R{리`�>Nw���{V���=^�!�^�*_���	�O(Qp�$u����R��X�'��0�`��L1�i������}�?�]��v�5Z�o-�닀�e����\�:�Y�A�t�fHj�4��cĒ��R�<���E6�)%9�qui�@_B���pH� �fb^�������kC�$��7I	����ur���\�UŅo�$4�����۷��?���2��]M��%�%�x��*2���='D~�0쁄:&+�����L�迶M���U3
�5#%6Fd�#���D��a��'��`����.���s쯑�������R+Z�J%S=�(�4���r
�#(����|��gH>jlj�K�^a���V��6�t���������������݃c k៶��b��S�j�̚d5W�Ӯ_Ԍ��C�5�� �=QQ���SS�����v�1s��J�^��>�%@�>O1q�½"���Q�b�@��u[ڲ*\e6ԁn������*o�1ș/א���9�zF�Ez��� q�%��+��K�^3������7^7A�:C�ۥ�A)��]�F�=����t���g/�S6�%��������ߔ� &�W%�Ѡ�#?���c�=pD���C#�< ����k��P:Vb�M�x�g�ͦ� n0<
�3��(�gU\��1_[���1��Ml�5vkb������k��O�}�6�V��وp$Q�PA���*c����D��@��(G�'��]�j�f��ru�^��Y�!�"�T���a�f2��&ީi�#�i'�+�ӗ������5�|�ůuu�&��<Al�H/�)���(���������wi<~:��#��"W�6��:=��1�M-.5��~��6��M�˫�ǔq�S�9�T�	�ǚYfRĹ9��@�9W4S��
��:�G��a
�`:��KS�B�AJ6�X�vs�G@��j��,��m*w��S�'(����!�&�rqKl��z�t�����X�U�3Q�LS)�q���&>��t�����$�nv`t)��;��^B�1�A��ܧܘ�.��J�/��E��l�X+'�A�pj�-�	���j)>֡��e~���ϩ\I��3N	�rU�xȜp�O&��Z���Zm�-�3�;����g�]�`��/G]����)Q��8!���O���r��nj�g�Y���r�`��=� ���6�����������|M�3'׆s��;1-��G��.����\;z����Lѓ�h��������t���N<k�|�0
��![�i4Tױ�Q�K�a+y�rL���z�zF�S�y��u��9z�t�Z�+�R��:#��}Cb�~?:���a�ٔV?͎��n�3�B�#P�q��c��+A��lb�;�e�5�h�#7`��ʈ�:�K)�ƣ����-��RhbA��?u3E�	wa_�|��Q�Eor۴�|�r�?߃�II	��l#p�`柨�m����鯼G�L��� �h4/�_<)���b��ޥ&���"�aZ����:�*�1��Aw��#B<nɬ�e���
�N��ɬ��H��e�@����s,���z#����;mc~�@��K��M�<�-c6�fh�3)u6m&�G�N��q���A����������)���+�iַ* 't<1r^u����E�c�2��M�9h'D/@/��'0�G��97�MopP�:;���~��M��r6nIÜ�~�w�6q���7=V;*?�����0ջm�_�D��:�:�Ő���õk����k꿖�"D���>LI�håz�R�<��adj|[����hr���5(4$�N�v�S�����r���(�6�������X"?�h��]Z��Kw�_���b;����	%�4�L+����HZ�3���~h�ˢp�M�Y��*Aq^��V`YM#����Vmu��p�K�#U�j�<v�'%�5{B��6��N��J��ư�J՗��{o�����Ϣ�EGxpl:I���Q�q�)���!�*�Ŵ�K�MV�TH\Sn�p7MP�v2��P�M,�[!ݧ6)Uۙ�C�R�{�Ӑ���#̙0�XH��9j>ץ7�@$�#i�N��~��h1 -+�%�B���PW���i�����I8� d�H�=.TJџ��,��nZ��	B)B_��2A��Q-�v"�o�w=�4X��������m�ox�VW6cH/�����D�N�� ae �U^��
����l�s�`M�&ŏ�V�v*�PY�dq���Z8n��	ɚ�f����{#F�뻖������8����x{��.�r�Xא���Sb��{��*��h����c)�Ϯ���"�~'+�J�M�=�>s��y<:���7򁨠r��;j�K rl�`a���Ku�C#�}�=���x�����m"q�V��Un,o�����l4�"e���/c�tHRY-��EXę�"�Ӷ/R���{�BTޥ�tL��s�m�)	�S�L�������I�_��t����p�)�$o4C&{vXE;.��xބ�)���"���!�>�$���"g�j����oo@�Z��C��9L�O�݆������"��PT�a��Ѡ�m��u3&5��P1�����]W��3�9�b��YOOR��� "������	�-k���!}���~rY;a3�������	-�^]T;o�$M�}���ؗ���Ga�|��NVՐ������]ш6��R�݃���*�i��M u�@���^�r�z��C'��â�x%9M�~&�	>.�U%����%>䤛�0乁��ޫ��'yV�;3�v}��<EG�+þ��t�����+�S#|���P�r����]w8�(^Po�\�	+ˣc<�>=p4Gđ)�:@�&��%��)���~�s���=)w���-�(�A,І9m��B �#�:��<�{1z���qr��k�a�����~�p����
S=��g��P��mrP	`�����m֍���ƣ��Z$&���o��j	bz�=+7����]�pO�0$
ZҶ8���YŷҰ�=)ػ�i�Tn�/67�g<��5V���\��,C�Ļ���$(�/<,����A?3���;8��3y�ǟ3�v{z1X�Tg���N�ןygkfO��U5A���^0�L������;b�/���C�A �Z$YU�MA�N����ԎG)H({BUikf�"KC���7����v�h_w�x�'�mҷ��GXWA4yan
8��f�{ukr���Tg��q	ن[ �sQ��/�pbH������a�,b�:�Sc�g�-�ua\;_K��O��E�1�N�7$�J�2^�:���;���O�P13��%�̼á� ��I
�~�02�Tm��3X�b^�S|1L�U�v��ZF�+L6�C�+.)"�WϬpUꚒ0� NYG-D��`�L&��0O��n�S+8^����:��qĖ{ز�,^�RWj�9��y�:�&��[��B��])0����Ɩ���	HDz��T�*2[0���[��Ⲷ�sl�O(�0�6TV{mz�x�!�b�9��Ww�W�v+��=���>kj� ��g��ۏK2�Z�E6[����sS
��G�ܸn�7�%>�V(�Ri�Y�����k�Ӏ�'p�2�M^��m������ؘ�����"nx�����ѻ�M��~\|�8�zk�����i���U"��q~Q3:�^��yww<�A������M�3���Wq��R��n���.�J�/0l�p��+�sT?����wv�}B��m{�?�-"�P�ae&��a0Y�b�mBv�C�(�R�-��2�
و0h<���4��Æ�
�����R�G���q�����I�7��m���D���h����f���0�7b�����8����e��	���*i"��) �|�ו5FY",�Km. 4Ħ��X;����r�\�2��㎟��w��{dB�W&#�|�Ƶ��ִ��cN�$��6u<W�x<llTLET��e�1���Ҷ�*KJ�����ΝK���;OY�5�Y��^��5)]. �{�|�(���%��c�`���Y�*��{���8�g9|���<��z��U��]:v���b o��FN4��╌&;�n�}�V
T�x�?WY�l:�&p����H�	�deE341�����6���ޠ��.�����$f�Aʊ�x���d^:���;;=Z�"$^�[,f�RJ����lS�Y���J,���s?J��38���J�88�4��k+Ipv4�����p�:�y�/'!�t���Qb��M��u�5�3����X��eg��N"�h������g��*�\�H}#���C�p,�VN�7j�{7F����-[�-��4���4,~�cwr޺#_��]�pk�hY�ҟs}��W����F���G���X���e��@(�e�nGʲ,U�l y��G���4��h^No�3?F���0/�'o2���4�<�Հ-��x�9��n�����k��Nl�4�����a�l���"K�:|w�d��Wi�Uk�5y��- v�N�ji��]�J��,���I�θ�ў�sh2�Q�����C��I�)I)Α�����-�>�xf��J D@������d��d]T01�R�_�M�B�a�ٳ����D|��Bh�_��*��]
Ö1S�⊘m*DgB$���)��6��o> =����Jjc� H�8�p/da)���iQ��o�-��v���N.[7I�48WƖy-����Nþ��[�w���BEN(����
A__>�V!L��H�u�7FK{n�����*Z����޽[��Eb�5��aI:Jߔ����n��b�a��X-v�9�Ϊ��T9����o�w�՞�E:pBࠦI��&N��>�bh�ΧX�M��>V$�q0*Z���4Wo��QD0�1�үtVlj+$7,?X-k�i�_�V�SbߧDS�߁��Qq�#I�$���t�4,Ĺ=A������0�隳k6�V���c)��t�,�P���eĆ!�Q:O �G�El��L�������}ZS�I��.1r�;k��m$��JHw���0 �:"#�������(݃�[�(��2�C���.6���(�υD��vY�\S�;����i.�?�+Ĭ�w���E4���@W�Zt��c/^E�yH�v�����g2<ƲŽ�u�\˫X��m�	:_Q��d̃�\��RkK������<��`���@���>������'�J���kd������a�Hq�f����B�^��9>�q&+/L�U�Ya��b��"#�wu�	���G��.��8�{�A�x�\,z*�#tȩ�}b��(n[�՘+�~7
����(��M�7�#��/�������<�:q��#��[���]��0�L<��������ghd�1�����"�9�J�=z�%���b���2����='��vzy@�HUy��;���;,q@�=�T����;�Tei��}p&��k5ߠxmU�2����t��<&:����=�
D�-��ʟ"e�ܿ����F�*�^�j��d�S�J�+�� sL�s��AM�1�LK1�[�X� �n���s���ME�H[#t�}z�G}�#ѷwl[����#>��ʃդ�x{ݏ�Tr<����}���5�~���|vvW7�?F7����}�(nSt��Wu�Q.�G���
<*P;�A�}$����(�c�h�����҄վ�b�j8%{��$x��2������MKq'�Y���3�X/�\�&"u�-���d�p�� �j��HBj��������h]����1k���Q6��h��_�.��/�$���S��&K�I�dI��^����J�r��)���`�aI]dM��]%�u�4�a���*FC��(x�*t�+9+�B�,��M���S�0�}�Oa3Z[�^U3@zK�Ӵ^D�
��㗈ܸ%�ڄ����&�a��:Tx��e����ũ?����=�< �%���E����zo�$3��$�����)?l�O���}}a�ɵ;2N�ѡV��0�q���G������{2��ǲp��1h�NW�GD��ڶ���+�h�>�������%}$o��&r�1���HCE��t��Nx3��,��Y:T�� ��b/];����>�����y8<��#�}P�{��h����E������$9��:VLaA����T�Vʫ�c�.��\ yta��n�T�Ad��y.<3{a�QP��}��e(��8T| _�̺�s���T3�{�<�T�I=ї�B�1���s��0�ӮI]n��*�	���3J���pS���`��a�o>��v&�6���
�}���i���rveIK�����ۏ�4!�q�oe�:�\��_LTO�Z-?b�
(Χ`߆ �U���fٚC�a���1d�Y魓���f��YJ���^��L�@f^6C�,���7����N�:1���K���P�]�ѝA1Ooxgl��G�2���x�Q��_�AkIED��7l�ER�z>e���Ga���HC�t��Ԇ���K�A��G������p�"�Q��u[�
�%����M�<���r���˘6[_��D|��Q�a��,f ���QT�Xr.k��D5�K��aC]�|�S�b���q�Y[�|mk:��M�{��I�h�-�i�D͚`k��3�'*��m�P%|�g		l�	bGs�>k��C���^�I��Ʌ�ᇂ�{є���	�F��4k���Q��T�3�]����n����Yw�lR#�9}�!7��-YO���АPs�3��@�0
`՗[6�=��%��ɥ�����&ͭb�d?�J��/gr���g]���{hs)��X���Y/T��r�bI�� �a��=�� �>����G�|�j�cl��mJZ@�Z�)|'�U�(�ode�H�m�:��<�-z[?ƞ�7�o����;���
cq,C���zJL��O����������P�g���\穖t+DR���b��1�_L����Q���DS"�����#"À.��rIt�,.��U�p1Ru>'��o����/�9UYj_"�T���1K9�<�v�f2�ꆨ`��Ë%��������=���VԌ7M��35 �Y2U���s}|#��3�,�O���|�!��9��{<�qa���g/���1þZ�k�N9��v�<xI�@[�*ȧ�t�e�r9��4���>�p�"��Gģ;h9jQD	��`�2K?N��㤢*�/h��������q' l*���g��bը�C� I��]-f�Tyb��	ޭ,xڶ��h���j��"(&��;!6�{}J͘�\Ϊ�}`^���=��G,�$� �Nr�,��m1W
2C(� d�M9������eW�������p.�`��\Rm��84ܴ��Ym��T��@��ŏ-�B�z�k�����q��\_�Cx*�['��:�ٲ���l�3�6~�g����e��|�Sk����1h�����v�w��ʖtZK�K�y;_�>�jޕ" ^�}'�_W/`W_�	P�;]�~�|���_F��=̋C�ԗ��Uꎐ?ᙂ��Hj'���_� �<�$+74��%!KQžW��¨��K�����8 �C��V�����"��@�t�L�r�s*��p7Y�E渁�(�8���N��"6m��=�\�|�'��z#���\���s��"�Ɛ�-����'��[����no슺�Y��]8���\�����S(�(�|�P�X��bͲ�cr�,����w�|k�D�N�\��$�m5qU�^����l+�Kn�Ry���}э7>B���>�^�>+i���t⒇8\�$�4��v���y�P�BE�,��BƁ�c����d���k#�%�FV9!���7V�˓�O�83��ߗ�,�,�ﶉFn�M�.����:+]!|J���׆�s�Vɢ��Ji
�� `��$�N-�D��h{Q����dϷu���j�̘�����\("H���{��`A�D��Å��V?W��f��������!�;cs[�+��7��GG����c�3��d�Q�.�zT�r���T1���=�C_\�v|8��"V�n�/��vg�Ɠ��ėL��4�)�(����k)�4����V��G����S�B��c1��d��v��� �ȼ�qaj�P]�J.N��x���p=	(���/����A�k������МM�+O��CZ���Y�.k5w�aW����_4���bt�/�Z%z��h'#>�o�;$,�}n$Z�v����Jw>�YJP����r��@p�]����X��5 �L_yT�/poþM�c���z�WD��:Vڞ1|n��,���� ��Wj�{��ԇ��d�t|Ȝ򇇼P�^)!G�z����33���,��Om߭;6㼖)h�\��/�U�̵�P��C�����,}l�{na[~Hhb�MnS�+�X]��O��F�@�Gr|��U$.�_2-����C���,l�$aZ�5FqNV��YN�đr��,��[,)/6u^��E6�t2nW��-rm�5�'���\s���ϙ�m�H��^�d�h�#*ʴ�]�WY��eJ���L�M��CA;�dm(�3�Da`@`���6K���dѶB)'#%N����T���X�"� 8j��)�<���4��. F�5�Yh����?�@�Ss�[���D�;�i5���ݶ�Y`�Dw�}G���r�X�G�=.��=�a<Y��4�Lʌf]!~;�Ǹ-NZ��V���v���h8�9����^����9e�e��t��g�)�E�UDVشO�!�P?#	&B�/+�ѡ�I�~�5�/�D�� �M�����k&�U�����_=ʉ0&C]�=ji��אQ�%z�U�1o/�ГBj9�
�&&�e�{�+�<�SI����鵌��.�~b	��Ŗ}�;89y2���p�q��۷|�:�ej��W�8e_TW�Gr�&�#�P��E��6���Ep%tl�bm���a=����B(	\�'1\���c����/����9a�b㘢B�cX��>�u�9ir�;�8������FՁ��)����4%`2aM㝶Nh�_=�������o#7ӺZ��uJ�ǡ��k4ԥ�d0G��-Dw�N�x3������#}����c�C�l횞�)�����K��H��a�����"�b�1q�Nl�JJ[kY���l��)'�uW_
�X�⧻c�7z�T�1��ES}��z��A�-��i�q�k��q��a9n����*�F��@��M��'c=��������N�-���2�HIR��[�h��<ǔ35�J���Sh;�l) �Ǒ:�l�m�\����p�EI/8�6(�6i��Y��w{f�O�a�8�ﯦ����u��Y�"��B�VY��z��w�gH:C�ŝ)\�w��.�����Nb��@�.6�}#���Հ�ɻeK�T cD�b���I5`����")�Ίg��HQ1�Ε�1��'������=�E���|/-����r"'��,�~�Pav���k��DX	�'{��Pa�+y�&� 9H���6�ڔA9;b�2RyQ�F����T�Y�g�i�kZ%��+͗����e�&P�x�jǐ:�%R4.���;Ql���])������s��fj~�n�p_��r�m��PB��i�3�0��p����a��@v��Õ���q�7+���K����O�g��d)2q!�2�R���8ǧR�}��z��{�<�!�@(R����t�s|�+q�A��Jb�|�Md�'X�����c
d���8s�n@�� �Y�P�I:���0����*�4��m�ِd��n�V���ܳ��j�����RVRkm�k}�w�Z�bc���{��NO��o	(�,���a�>P�1�#���x��~L�mOY��U.�%P�}ﻣ&q6��L��B�0��{D�TK-_(u`mzx�����ko���M�کO���_��r�R�^Zԥh��4����u�G�Z���{\�����!��(1��FHI�
ʩ��(����|��W�@��16�,őT���_ ��d]��#_�v'��xl	CU+KB1� �Rg1mB�Hú������������1N�c?�� �?� ���G�U�W�Ʊ%9p|W�"�)>0/�{N�}$�YG�����z0��S���̼���&�=6�)c~�l�N���,[\��P����J&����l�~i74R�K���,q�+�I�/�N�2��e9F�T������P��s�$@� +l8N6.���Y��?n��	U�V�	����Ȣ;B�k������WÕ��n��QA��}3/k�����%?HX��xI�� [te7i��B��B*i�X��(�Y2�,�8V�]l�,�x�� ���۱^��f5܆����}���0��?X!؛B�_}���*-^I�7M���vP�P+H��;���i9R/��Hy�F���ַ `�~	�y5�"�u�)�h�#����}	vmIr��_JB8,�梢[9�H���wy8,I$hg��؆�%���0!��t�ܯ0�蘢 k�B�)H�����[�?�R�Ƚ����[ Dpe�ў�_������&�{
PzYE�������L� �R���*s�����u��}l�ܼ��	��s@Ϙ�Ӧ��t?���`��A3 �����hQ�,|*C��:U�%���;9�����d�$������{lh�2BՈ^���w�.�I�
��進;�99t��!�viZ�r��/}0ԛ�xœk�e.�p75$S��<���N^�
������X���v��9+<�[��͂�%�f�4�v�m�
l�0*�A_���"_�~EF�Z5ެ`�L��Ԯr��fg&�܍�D$�1�n�/9g�2�sYG���j������xX��ST^~o���'?�N㍴�d`r��B&��~�$�>Ce����5�w^�����E��^�\J�7c��]7�<����F�{#O�*����.]Cpz\]��x�*��!�[�����FEzb�Ǩ�Y����Ũr,���k���7nX�}IMx��U.U����[�K- �D�ٟ���8�.z�������
���6��3>�[���tP1� �5��1�}����a,���`Lq����kz��ڲ;�y���dˬwZrc����s����d�5[[��_-�9�o���o�A����N�,l����Ȅ$��n�6?��ݷC��vKg,4p�Sе�ݢC[</�C~��AU�jT�ȸ���m*�����^}�u��D��9�}� 9��(I�����1!���e�,��0���.��Y����MI�(K�iM�d0w��u��=�s,� �e�&�a�ê*�4R���c
��hK���׸�A�D�@v.=.bƯ�CSݣ���_g:#�<�_�ʱ���|M�^��IW�dq�2��0,���J=���:�kT�<�0��Zp�����׃CU*d������e��p��ԥ��뜞�`&�p��E�d��o�5��xȅk|D�S3,�_gi3�3�nqn�2�<P�cPb�?b������xM$�/���*WE˝W���+=�'��Y�Q)>�k�ק�=)�i�9>G$�e�#��v�W�\�oJ8��ѵ"e�S}w^d�3�]-nW�^{24���۝�oy������q�Q������kc�~�&FnZ��OYPz�����m�%ߌ*���/ˍ'R��?�B��H�O��2l�O�E��$��H�(b���=�̯	N,��6�x�R_�&�2����V1��
�>�c54�Q�HS���6y�H3l��vJ���d���O�L�Pk��x�6�b5�`&���.�o�4fjҞ	/�X����g2�'�4���;�d�i���=��yn�r+|��7~q��5s����F��~�UVep��Ϧ���6�5������p���--W|��3|g�R���5\Vp�,�}��J���㘊��&��6�I\e�h������9�ӧ�q��`���;�x�Ԕ�)e� g&&
�"�X�"��)�(��Wyr4��i��*]l=�f*�F�U]d��ʖ����4��3��U�Z�.����E���;�""��|4ò<XlA˪D�����s*Ai.d&�=��*c�ѵ$3�YG���ZP���=��E����	�h�6%)6Ys��nN��a��)� Sx��p�`'��'���{t	�8�����LCdX�[Y���i����%�&ȿ#)�B�lx?��d�)Ri�;�L^!�!��ޏ��n2:���{Ȼ���P�E���-��h��D��~�%!h��Q��L���nL�b�69i�G���9Õ8�9��D�0m.��1� ��DQ($�;��,�而f�D��1�7��9�N�[�N*$�_���z�Y��+qc{�Y6�uR���-n��X��C�ǽ,*\Jk���>5d�׉���y<�
�ܗ((��V�%��]�@�vA�����a��rBjT;-^
"@:�-��/�~	��/�O������#<b�]zZ�عՕK�\2&�]s6�)�2�y5��Ke���1�;������-X�Fl���D��|.�,{�l('!�8}N�w䀢�����Ry߉FP��Z�:.d���)[���k�m�J��db .t<&�7$u#����$�51�U��0FDfDX�3��߼�+���	d-�?��AWr%����\$�es�zT�&��Nt�~����d(��#l��� �􆳑�@{ǘ����;6�U��MB#�Q�>�>��4�Ʃ�M��������l����'.�{��X�����u��e97��͍R� ����3_��)(�CPnVp�����*7[�p��&��K	$���	��M�f24#��'
,#�r����~�ڸ]�)���4/��u�J�k7J7�N�o)}F���qLA�kf@r����dP���R0;�)lo����F�<���¹�2�$�O}�S`l�B�*P~����d��������g�Ѝ&r{�!S�����������S�ڎ�UN b
t���x�b���ìe<�/����b��#($��-��5��a�H�-�����}O�L
�^��H�l�	b��m��"߀��:���
�8��')�5e8��-�z5B��Q#�?��Y��̃@��f��gs�ի�؛�ٱM�4ͳ���͆k��k� ��s�S�����H=��\��MBI�t�2�����K8[�����׮?E���q�����6P#)�@��s�FĆ��p����g��0�Ƃ���v���{����^.��կy�;�%H�B����@�Yu�$yFb*r9�O�,�������8�6��#@k\�](δfs(�v�/���xM�U6���;��^.hb��6o;������u4������^G-Z_�-gQf2��g�������H���lOS��C���(�c��
�S���,���Â�!4��=��F��p�� ����|kv�
L~N�<�#�3����j}4�9���C��&�f��tk�tE�%W����Q| �;BޣnЦ!�A��h⚈y�����Jů��@�'r��T�yz5l����K�Tź��\_s8��j�-rTΤ�1���\0p�GK����y�EM�����
�G�Z�+ �)M�ڛ�!�|{��{���Om�C��3��fC�HF�pVViBʤ�h�T 0��
n���:�|J��g2��3�ʺ�1Ux�uf�L��i��x��QzGU���
h�@[ٿ@S9﫫�_�M� �!���$�8n!⑰��Op�!z8�b��a�D�|��svT�g�HC��;��+�2굳���5�~��+���)g H\�_'8<K��E����=�\Bb����*�q��Oy͸U*�Y��9&4�T��,���{���z�߈*BG[ݍS=�#9��p��YI���*&�y?d��U��s�c"�G�]{�{���ȉ�1�{��w"ޤJ��e7�bY��bu@��IVE�*��:�O���
����g"YZP�_6(���:�B	� ����nc��}�k��_V�L�~�z�GS��R, W͂[��;���0MΪ�A�XA��iFSΝl��)oD;V}Ao�@fɮ�%��Z%!������c}��G[��\�3Y�2.��G8!����42� Y���A���lC��R@��A} ��x�l@G��;"8 �`_9��m6�[S���:������/+4�K�O7ip6�G�rE_����������u���A�� UH�o#ֶ�]p���E���
3,	;�-4W��Y�U�5��V�S2�jm�ƌ �Oc%b����;��C%9������ω��\3��?�֚Ʋ��F^��Y���W�74��Ǽﭿ��(
� ��ir�Sç�D�S�bgE�����Ͱ{��`5:�������uH�7�7C��5d*�zG�E���2}0�>��C<�Ol��(���8Y�}��(����Cq�H�K�ϧƵg�{��A�Ud����^;�"Pj<@����F(p��B۳(�DE�-��l@�v�;���N�ŬXm}��|H�?�d���p�<j�LM�yo3��LgTH��s��֛��1&� �;�y���RN�L**f�wn�� ��l<D��G�2>U�SU��D�O�H�)�0&��[4�4�����CEv��[�@r��&�-7���&�;~rM�,EZK�@%�n��ł�M���/v��ƕ�m�A���A�P�w�T�����[?��Z!��|����@�i�,ծ��o"�T��,r5��R�.�����Ѵ*(�$wQ����S�5bE{�7�g�Hh�t����GBa(\��n��������%:6R�w��Z*�Z��Ċ�
Lh#0D�N�Ei �!�AJ���n'���MJ�T;�2�5���I���Wr�%F��\D��/���hFD�3*pf����V��I��jg㥠�I�ۗ�6�!�N����󊑂)l��+B/P�����=�;�Bfް�$�4)��.\|lU�+toe+
��.��{��]u����;.�*�G�z>��|?x�,J�To?�c_���R��2������jrp:��#X�ډ�.����n{�ǩ�8ɽ��׈��p�?Ͷc�~^ݣ�(�����9��e)��$wH~�(k�×����������F2�ڪ6�	��ze�*����{�پ�n�5��y�bL�`��qYJ�?Qn|��2λ�Z�x�A�x�8�K�]�ð����l���%��Wn��J�̶����ľ,gw�ˢ*���a ����(�ϙ[��2����"���v�|��Z�gN���������2���-����r���b��~�Ы_a{�:ZIk���Fܞ�@Xu텗r��ڻ,_�P��p�����[Z���Bޖ�?�B�X˺�ܙ��ޝ�d������/
���#�����@)�^3��1[Q5�Z�'�0��^;�%���{fΚ�W(��LtR.�s�S���s��H�����_���L��?�q��o���Z���3�'����xE~D�k΍,�'b*�K,C���va���N�iz��'����I����^5�$u0M�g?���lS����H���+H*���f��s�26��"�n��p@����F�U�w�2K��a�fr�rDY���	��,|�j ��J"���g�3B �&�5�<�l՛��BKc�a��� ��Z;\8-�.��1�X|� ���]���4Z������w�{͔[�K}8��O�Sn][5�;��.�q��K	��3��A�|4`��pX
�jҪ��{B�e��o���7MdQ��w�^u�����|%��a0���� ���\{�+_�A�O^�~Í��x�9��3S��i�V�X��r��uPQ}��#�J�N_���h�r��
����S�����EnjO\p�"�u;`���]�P����9�����%��6�v�_�=�Z��p-[��VQ�-L�����SK�{e�˿���.Z"u73�Nd�js�����.��!p��u�r�3��_��Iր�`��猲p�w/��n���(+�2 �z��q }���x��5��y��e�3���ݻ����
|&�uQ�Mz���"K��BJ������7���qs/h��e.�m���H�:'pS�����aᡆ��&@���vv�2���"Q1�Τ�XN�+ҹ���4�k��i��R�6�p@�2bv�i��~��4r��1pz�O�p��jy�����e����CkQ�9�NbԘ��V;Wfk[�G�\���>1��ʽ���GC��L>]����,�Z��7z�4���	��>�ѫ̹�䟸�$��zMi���|��8�2�m�ƙ�)w���`��Km��4�;zB��F?�p��!��f�NB��HKZYŘ�>c=:^�R��X�b�5��<��Q��r���lX��0���|:e[e�K�:����N�[V��r=��h�A�r���J+8����s����<�<v���a��wbK��,T7��S�/'!,z�t _��+b������3%�G ���L������T�o�I�� ^���<�#�aȸ�b8	ͧ�;�z���^F%18�ӷ+�:l{�?�뎏&7�(����������{uX�>�C������]�`��W�]��ư���9������!IRe���pJ�WV���%���[Y��B� 6(�F44E����$\W��.��~�$؝���� -̡�~�s�n�m.莾`]���h�l��/���7��&@a�:��(F��2�4�x"��/�4.��G�h9�`ט�.d&�W�� w��/If�2y��˫�B���n�,
������Y�����ݏJƳ����24g�!�0��46��]�`��G��v�E
as��r����K��o�E*�I��x���FJI��4���]s Ѿo���7����I�=[iW� ֱ���=x�,E���@j�R�h��N����ßs!��ӱ��[�y�5���bMڞR{3����(�7����X���:d-\G5D�I�:����n���!D:- �$���3I۵ijҲ��|t%��c<3�<u%	%���y���� �Lw$�VF�=�WV���L���o�iW�>Q�����V��Vx��
��5�	)eE-�����q�����-� ϶L��j��#[D�2='�=�}U'^y*O�_m�\�A-8��,�3�.�Y��ĪQ���H����j9��s�6X�[
c�
�
e����Q��&��R�?ү�h�F.L�����oi��*�C�E�'0n.@3��	�R�mr��C���h��q���I����!ip������0�]2\
�~+&z#���+�)Q�X��2)kfw�\���uǽ?IB� ;��dG���w��Jc��ֽG#ǭ6>��@���b����Tup�2�|x~Fc��Ǜ!�F����dQ�GJ��6��)I��a�NT5Q>�AO}���y_�����v	?/�Bx�ʑ��
n[kJ�ё�T?�Wgv�����J��A�~ix��1^3�!K�N����2���.��Or�ϯL��;^mZ@֡��@T��,��U�����Ҿ̹��D%��0������w����L�raҟ���A�1&�	rK z5��^��j[<����prx &G�[��e���D~,A�J�񽪒8���LZ�̗��+bT^d�-�L����|���/HCr\\:
��7ڳ�E�
qv�j�=�e�k��Ms���OM�I�B���,�2����n��h�w{j%�#�[A�Ⱥű�Dˮ&��9���l9��g�}v4[�~H�f�ջ9pz�)H�s��[�Ja�d�"���D:��f�r�t��"��KE��s�Pt�~�O��k&����c��R��� E|�.��祟��{����跾I.�pa��v��)�e{�j}�cJ��H�́N���!{��ȯ���|��N�J�-��le �ދ����&*�h:�*�'��$7͇�ς"݃���X5���F�U���q�"�Yg�W���gP.�[�{�lU0K&=�hv�2��!�:���`�'��
�=�ó?��FM����#׽���E���#ӵ�\�|t,���(Gb�rk�o��a�� 싟�"�>dV철�-��׮x�D��O�0���(�u��.N��
c'��˞��z���6�[��=���Р�-B����_ ���/��)��6���t��E�SPD|��������5�Q���q,��f>o�5�N��0!ߏ��x��,,E[�%KNr��&iPq�~��U� ����g l��x�ȯ�{Ϯ��5��̰�V=PֻOo�ʬ��w�P[b?�0��0t�R�V^�����RF��Fzl���繚Ҫ'c�^�қ���\���������S�(�|�c��}���X����<���'������eB-B����xU��Dǜ��X�ΐcE� zڤ�ko����6�E@��f�iH������6��
Ͽ
��2�Ҵ7���F�^z��te�]��R�O��u��dO9G���
����ג��*|������8�خ<li�W���)8oR؄���fj�o?����4��SB$��ָu�+Ǩ �1{�����X�՘�����`���1'-P	!��:��y�XK��v�Cb��/]Hs��&���)��T�`�?G���+��c�d�>���[�B|-T����F�E������u"����My�t��$4���t%�$��|��Zcb�*���⍞3��W�n�y��)>�Q�%�51f���ў(������?D������V���T����~�>C�D�%�6�M-m7/l���H��^���%DKE��Ѳ��[$Xp���b�l65T*����BG�ԍ�Xw�O��b@��cI8kI��׋�X�lB��g�U���	Ч���&����*X���������-�ơ�����"�۞Z�OZ8lѓ�ԛ�bF��Xt�b�<5�. �S�E˾�'Xƪ��h}���Ӷ��]	w�����}��f��f�#�3[���dU���6�:�3F6�G����`[�Q��)&�ݓ�n(��OņQ� <̵4�N4�me�E�	��;td����
#�Dɢ��o����Y;9�l>*�"���A; 	ӕ�����(���잰D���91,�z�{BY3j����u��E�G��T>���s�G`��G<�d�`�)mt=�@�:,�؆�����`oFr�����-#Y3P�x���@��d�y��7Գ<�Wr,�r�`VF���z�su�r�r$Մ���ӗ.���r0�])��Qv/=���������P��zA�=~I~�]D�@Lޕ�e��4}�L	 z�E�@u<�K����T�Zjy�'&ͯ���p�����ci�]=H�m����xF'��b�i��ʀw�eG�{WI�о�E�s��>k&�3҃����+RԔ�6Q	ZK7dLN�W;��%wM�žoQ��"j�b�D�k����[E���?�\]-iI0�=w�썾��+9�����0�]$Ĕ�\A~a�р�aާL����'$�4�����w¶��{$���q�$�g��j����T'gs_�"^p(/ݘ���8�ƒ�MX8���pr�/���csFC�;V�"4��L`�~Wn��Z���5P�)o��`kR�+� A���[��bJ��?����K�P�2]"�WM�>�H}{՝������ U��p0_�!?̧�f���"����H�8��)#�b�.shNg�~����5ס;,��I`a�Jϕqo�E�jj�<ϯ��;K@%�
^�/($��*���J��������Ug�`��� ������3"���e����W�!r��=0���"t� �~���&�;!S{���*��aA�J��6{,�a<�(}������=�s:��M�1V���h�^�����ՔވF�3J7S�Ԟ�*P��xrH�P�)M�'��ᅰO���Q���b$�cQ�DN�n� "�D�ó�-�8���b6���2��UY��0P�$��>��/�3�>�,��E�)�Դs�V�V��;�Wjw����	zG����>���e�+~#���W����_�@�Uu�_����Ë�����L��
e�~Q>��&ȽeGk��Q�aAbp	�&n�g�0ŀ9pPu��áW%�;���@�j��{Y�I�;Q�����������y�x�@x:�5��JdL��b	-�'����/�P��,���_b⨁�ȸb�U1H�k�s���E�C��v?t� ����7CXw;yE�~�%|�
��֌)(I�h�������8�>YsSg��^5���:� ^ټ������F��@βi�T
��[�_�baC�l�D䜪'����V驲�қ�_��^�ȑ����j��	�Ҹ-Q�p{7����ffg|���7��
��c"�F��'^{>�'��}>���]S~�^0w�5��}G�E8_vgK{S6���mۙ�B����y�h�u�m�CLN �[�t^À�ݐ<�������%(�"	�h���i���^S�<��04�)��?:���g}`e���F�~����adhj%X��v$S��/��(�����.Rq�4�n?��v;��O�Է���z�SlP�g�\�	����#Q�Xe��%�dy�@E����Dl��;^�R�p�pR�*��0T1ܰ�z�w�_�T_��zw����5�����z�݉+��H�֤/)�A�xO���k�k�c���m_+��r��!Nl7j�C�ȡl���]��y���>���&����Њ�qz�f��D��^���M��4oi>������5њ8H�(a�"8*>rGq�jH�9y�Kzp�������g.�^��|��_E�{�,�*�g>�(pΆτ2�tV�NuIº���QW�b����d�ჿ�q<���������SW��c�pY+&_7�,��W/6�;E�!�|@���?�6�H#��DVh����ڶ�g�V	c-\��[�3'���g�iF�ļ'g�{��Y �s��>H��jz��?��q�	S>�}n�������d� !�;�T�݋}E�f?�M��P�f�h)a���r)Ծ���T5�H;���sϢ�o�
�u���UZ)���**�݀Ew13Cf��\Rǉ�;fE����ݱ�����i�y�2~��OD���]������m���{.'e��У΍_�9���%�}���Y�=/ʵFc=���Uj�'���n��Ž��	����X�$�{H��۾�F�E�
>�Z~�����W��ѐ������$�0:K�rc����d(�Pr�W�[_���
'�W��b����Kw�b��+蕅!��Q�9��BE�	�2ط��3ψe|A^�\=e��\���q�a�s(��q3w8��6�Nk%�=�=6�z�7U��iy�$�-3XZaLƚ����Ll]�Ui���L����f�'��v�=�?�'c�Ս����bQk��_��.��b����qQc��1�X�<�Xk��lw������p��	����%��,���Hal9S�������I��=	��&:y���!U�Pρ��q��{�+~��N�:����9xI�ɶ�6"u�U���o$�$=�E29&��+���4����Oޥ��`z:6��<�C ?݉m����f>�V�
hˈ'}���7r�.$h��\@i���>�
��LكB���o�ʡT�Q�i���W~��d'i�e�I��Uץ�QP �X��7�aV�#�i���_X��*W��xaQx<Xo+��<�i���"59��y�S��$��&�^U��B��+��E�+�I�{�'_I��I�^��-3�_l:S�I��'Kf��gPى�D91Z=�����,L��q��/hЉts�����J�`,X��H�	f�x�,]�M����vi/�@����%J��[k޸߻����(��1�6�` wc���oq���AގƮ���Uｦ��A'Np$a5��lЦ�5�+k�@��_�/1�)�4ǢJ�̴�R恻��儰�z�
e��6}1����c{g���J����x8ȫ�hL]�$���!vh����S��F���a��*�GNxh~S8�;�I�y�\��Qz1xԁ�p\p����L�f�q�%�AGٶ����~�+�j�ʪ!��J-�(:��]�ݏ(�-ז��)7c<{p�����8>�ZUk�~q@�2��h��RUC̎�aұ�.о�����?�B5q���?@�Q��m�W\���C.r��9�I����җq�!�`���)���������}N�)WH�s�G�{Y��4�핫��6�U-�5����f�j�9�`%f7'6dў����]I�3��~�?��R"�C�4� �z���U�;�B��y�|��2�ɏ)=/#K~����yx����cR6w��1{I�wE��	>M��9v�����@v��햞��bܯ\'~�s<��@6x�N$�O��~nq�I㰄�i��z�q�-�����Z��!��{�N6�e۸Q�Ԓ�a�	�{?AݭR��v�v!%kݻ�8쭙�'���N�-��+}�ۓnOB�E�C-j��9|q�&#�<{�T�W���t*M��.!&O���i��da����m���(�<%����Ki��c�쮵�~�.�
PBh]7���Lp��@8�Pܻo�_�)�ު� �B~Ɗ�	`h~��˨�FI@�+gCIj��^��xS�������7�M�}3����_a#���?c�]����}.�քk�-b볈b�ڙ������<D$���niQnvɍ�[ؓ-L  I��\��4������rf@�\��o�2��c�Z9eaka��!��Sd]�S�V�V�
��>;4Vg;�[)��|����}�q��8�i���, a��r�W ���L靀�hL���0�w�S��{�XД�����W�?5���w(\8�����f��z��YN<�n�@�46׼��7���;c�5YL��k�a����
��|���c?�*�A�Fn;��8Q,ɵ��~@؂�Q�E�N!��x�>��6����'!Px�]�#yc��Ͱ���{D��t��Q;��HR��͸bW;ǿP�<���:I츭.��`�KB3¹�~��5D���G��>�5�Ρߧ/��������'8�=�6�mW�Y��2R=�taA�����f���O��@�k3���銤eZb{L8\�~x^��{ukt�O� ȭ�Nٜ��G�gD�ϳo�f`�SLPe�l�B��s�oOOg��o�?�[q��V�d��.������+��D�~rI��l��;j:t1C������Xv5�.H��q�.g���;�䆵��5���ϻk�{D�����g� ݏ�����#�>���po���<�dqi�lN7��g~�v����F|�f/Rb�ij��Un �qE�[ToxاSI�>�|ʮ�f��Y���n>�4�I3B5W =��� �E/d�������"g� ?'	�@����X���_�*\s%�����N\��e��J�.��-���xg6$!�&���Ѵ�v����D���՗O|��k�_���X����S�� ^�U�fd1h� ��r9]�K��`j�t���t�)D�S������U��
%Ǻ�$��)$��GGX^���kxv���'���#TI��\]��q��@��GY�(f�_=n[�FQ���N��JV�Z�1�{��L�o�w�B�E�X�n�����a��\ৈ��g�y�}/�=S	�#����< z��ު���h���#�T���V�,"|�o�1�̂�Ί�M	�p��`��*�w������|�u��B�Rl�f���<���`�!�3�'SV��� �gm�SE����aYl�p��%NqZ�o">��V�>؃�������LP��叹�qa��R��Q{=�O~f�E-��8�T����D�d��<�$d���\��3�K���	��N���O��Ǌ���xA��RJ���e6��N�~�#}*��\P(�v�Č��F����˚�'�F�KR�o@��L+��}��ԛĚ�U��\��-�N*\���$W���$<�U��<�:�\j���gR7��T��C3t*)W��tNH�E��y�2zae���Ľ����1����c��8��F�o�]�ce��ֈ�T@�:�wT[6,�p��fC>����[�����P)%2�W�)���F�!hN��>{�
�yZ���&N�Ty��"��kRgQ,����E��k�z��uw/[�4i�Tƛ�ZO>���'�Զg���h�nq�o$�G�����n��$8��V8pd�ϣ�e?ȏ����,�H-�����]l�O8�eV�V���]���3�A%p/߫	:���:��Kk�����Uov�M.E�N�q}�j�"�yǳ�ń����'���O��!M�H9���iܶH�9�}Ru����+0cyuТ���bͳ��ۂ���Xm:[��bw�q���K�F��I�,xi�%����
mOo����H�A��߂��ZA�����ӊ����b�:��e9��ߖA����3���Y�Uj�J y�n6��G\p���$�U�g��ޮ�{�����%ě�e�S����GF AZm��h���B��P�}�Zآ3��V�DN��R�A\�7�[���=�y%Jj�4��;g�,�?��"Ң� A[�ַ#	͝*]���v5��F�(�$�@ Y�A���EK�]Z��gL{�m��.�:*�	Ĳ�ve�$Pb��^���QymӪɤ*<"���m�ǁ��o9��u�hrx�Kk�v����"����(k��0��i˪a�� �'�*��D6)U�D�b����z3ܿ�X�w��
�D��/�Y Q�"����1�B�k��CH�
Q���U�4/��� �� l�JJͣ:C8�����W��K���  �h �ώ�R$��EP6�o
���`�w��v �R��W5�@���(M�n���akn�23���l5��W��Ti��I�e��߯z�sjf�ؒ��s����G/a6�~�'�����Ū���d����R	����-�	ME�d�V3Y��\E�/韹�ye��4q�{�f�L��7��m�@��V�`�z!�kI�ək���ۢS����p4�u���h�%��{i�rb��ۄ]�lD�1�2����x����h�Kb���R����I2	
k���<��Uye���D� L����q�7����4��3�/��x?���ϛ擥	���g��O�|����$J;6�'�4� �E��_�祩�Q�!�D����FH8�������`?�'�
i$����U�*h��b��MH��`�D�۽M����Wr*�dDA��>[�z(�.��h�K���p<_�����Y^��@b� \��:Mo��d�i��|����.����٧L�_ݨ+Ǻt��iv5�ٳ'���p��'���;x���K�)T���#F���JCU�ŭV�ĉ\d�A��
��_b�^F�yi�l��>��GMf"����9��uF �< -m��Tg����ͲX�fD��	r�-%C]��T�����mP�b�\ ��F��iu��ߋSc�Q�+��)qG&Fu
�+^��_and8��6���ۻU�d�a���Z���;s-J �E����J9>@��MSR"�즻Kp7\(�q�R2��r�eL�`�����֌5d�b���+�q��(wL��a�M�[W&�#�� WcU�Oט�U--A�&(ы���fX��^O'�^*L��b7㔴�ܱ�LJ�x���s�ןк�I�_I�Y�_����ɔ
Ŋ��d��b�Q��F�Ut�E�jlDP�ZUm������F7O�2f����#����`�(/�{B�Ne�Q�r��������Nj��$N�f��孧=��]�F�_�H�#����T-y��'E�o|�q=l���!j��MꚀ���H��3r]�~˃��� �p�� ��n'?)�M� 	W�ڗ��"���N�8\�>0���Io�=�s�j�*cݐO����Tf����_��Q�>��K�U��C�[3*�t�j\�``��{�x�x@�Q�qP�h����f����b!ѣV&��)`��5�ָ/�ZB�7�wd�Wԍ�T��SA��o�y��k��9C1T}�lR	�",��^I��#z���:u]��̭�&C�b���2���kS�{��02"�i@�4��&���)���Zy�(�+^�Ү�U��sXN� -c�K|Ffנ�{N�P5�GW���Yy��!�K��&��.�U�W�'��+�����ex��ܝ<�<�;�c�@-��m�B;�9("�h,�S�Z�e�ŭ�� �v_���:��(K�'��"4��L�PEt|�,'s�l��~���d�I�aХL��D�^>&�ob�������w ¿��D��F$pe�͔���
���B���U�{<g*ħ\�٭��ն��d� ��6��)*���_�t�&��51��"�I�K��]J�?��-n��#������r�p�1[�G;8�7��������	y�2�(��97���:��5;�_��'e)��m,X�K	����&m�-�4U�E�YpS�1��N��*��w�Ơ(�^VR�}1��տ���av�e��d��/\��Z��+�e� ��`j�d(*�Y�NJ%��W��ĊKR�F�E�c�*�H�M��0��~A�q�'-���7����TN�Tgۀ���t�L8��E,G�A߳��	Nˆ�tu��=�ݶZ�&L����؟��[!0�A�� #��!��z����k%IU�{ƊIH�@�I"��zF�/lX^�{N�)ͣ�RL����zj^�i�e�y��
Ϭ�?�:nm#KJ	�C�j5�hӋa���s��f^̯�K=�����hw���sI�Ds���*�X�R���ð����� ��\�Ihp�N1&����Aʁ�Kn��R�2���Ew�[�w���i�.��`}�����ze�a��X*�h�4լk�h�� �:����@�.�
�W��������	�X6���J�������<�/:�NE�v��4��� �"Ɋ������~�)_>V����/~3 0���avn�n�
�d`\_l��v5G�]�1��8�3�2{�`%�/��w�%����Zũ�� ��e�H��Ӻ�v�S���~��	�Ԡ���{���vݎ&�&'<w�v��<��5��>�v?;�+�T�|���B_���8�����&{|DOtȜ�����a1�"Q�QNoBP²}`RI1�=J 8׵�#'2���d�&�JH�.���)Bm�(,�c��x�}�O	����������ۤ0����w�+� ��^[K}���֋��D���Y/0Lt7<']"Q�-+�N�����ZW�կ	�&2�T�c�z��ˉ�w͓Z4�%3j�8�5P�J�'��� 6�*~�;nX�G���Ra�zE��#��ﺤ�(�0�c|�n؉��t����ٹi�jn#=D$�S>��Pam��e��V��\��{��s��VQN� �H�re���͇_�$��̻�A��> Ԅ+'*s�w�c�`U"7>J�"b������GC�L�׬�����z0�DǡrX��#��ݙ���,�m���}�H�6L~�$�H��E�9Ű�G�� ���}D�?J�<�yO|�5���?�Q�U"���s�F���N5v�ӱῇЈ��D+r�*�t�dp���*�eu�G�"37����J�DNo�kY,�v������!��O���N<t$?��D��dX7��#������w�I�f�rd6���>vb��^�J������w�U���Ag���l;�27�B�\�@5���u���u�`fca�ySI3��[�,N�v!�@�k<0�{��|၀Yגw��s�����"�p�5s�ˁ���w�:�s�B��*�.z\�5���olό��ޝ��C!�]��-�f�Z�eS��}��8�j��79�l1��a�y�M�P��Ƀ� Po��L>��9I��7�
<�N�jPUL����� �Zm��$>����e���S����T������0a�M$f����EIH?Va��;Gw�R�z���Y��2ƭZX5��5���z�f��7�٫�f������'�\�G�aDIE�桼N6��
U�s8x�)��Tv�]��CU�� �js]�Q=7Cpx��؈����9��ˣL�=Ù>nH!F��c�=&�m���@��'�dx�+�k4�� ���d6�m_f�{1J��a�"�=o$����\��H2���M��\���m���.˓s�'x��:Sz�({�����eN5#�=S[�������Q,����:�����4�:�0�s��] ��2�I���򐏈O���.����6u�Sޫ��yh��v4��G0B4E�'ԼK���9�vSṕ }(0�}!�ip��sX��]�q��Ui��L�.��**0�^���kx�R�IF��Bd�pZہ�q��@���siJJ��2]��_{�E�:����F�M��̩��!I�9��[jv���P׶n{�u��s6JU��C��^P?����n 7�q�����n���Ϩ-�޼���;K�W�i�Z=�؉y�P�w�����nǭ$YL���������͉��±{k��
�@�6�᥼�U̞�F��寐� ���p�𾳵�#[��G�So%Q�J&^�x���`�cF��2��Ȩ>+��'��4qVaD�	J������Z�Q�M�Χ�]�л8'����`�(-T@)k+�.�)�3���^~�ĥ�����B2[����N4��R�̕���JsF�V%1�������f����KG|��,F�nP�����K���+��@eI6�MQJ8�TJ�nb����%�@5k�E��[	���݊�I@G�j��dtT�@au���V��%�lHm�
���!�;�L�����O%�Hsr%��m�4f��/��<P�a�`Wר;���DԮI��o��n� ��r��!�D�V�K�H��N��~#�Gt�7��\՝�bHF=P=�r�5�6K�&�H3�ƛ��q`,Dɺ)^"b�13��M���b5��w������t��k����..���ق���2� }��Yf��~������=�}��Lh��wɤwos���ߍÞ�_B6#�!c8,�f�>� �c��Z)�|V�Ly�q;p���Պ81H
1��re��]m����=�0'yAMHt�1�=+��ʮ~�յ������ܬ�wF��gm1⠔a�q0p��=֖H Wt~����l�����eG}e]��H�^��g��i�˥k���pu��\DpۿY�H�6�m-%`3��F��_Dދfz��*]� �&K9pU2C����m�2�}�@�2�'E���^�xU�ꮷ9�a���vQ�`{�O��R7����\�?۵M� �������HJ�Qz�6޵��;�A%w��lRJ��H5�U¥���ey\���es�V(:�8�#�%� ��s��+�nz�kp�N��ɥ�{���o�C��\4l�j�z�'[\���"�QV���NF�������2�KB���A�}����!��~��JdoU��O�E%	�f��7�Dˈ�7v��PH�~�`���ө���,���G��
k��`;O�Wr���������x�*-�f`Ʈ��SFUy���^6A�X�~�"����b�Q.G0�#4 A[����2�	��N-�V� S;�s�l�qL��~m�ڂrPCs�Y@�$����5�rn>�L��[T�:>��K�;-!��|}����%β6^pr�:_ �ʝ?ݩs4	K,�+�v�E����#��x�|��P�����+�E$��/���S��u��I�C��c��T�6�HZvI�9��@�L�������I�ץ�g@Y�����ù�Y_�9���P���-�1�����h� 3�HV����?�I[���&Rw�^'�xi�L�<?XŅ��oX��7��Kv���
���ӟ��j�ٚCg��]J�h�����\�O����|�!˴�"����x"���
��B���n!<n�(��#�{���kW�+���᩿�C8��>'0hx��@�	a�2����iȉq���hr��h~�����e�ieEz<@�!�$���9C��K�z�H�i�e�`�{������!�4���ڠUԮ{��R�pca46ݦ���{���E��q��i4�8�Ѕ�ͳϚJN+�>!��;Ru�=b�o/�4���O�],���y7𺦎\|�2K�ocSOJ#[�R�u1��g�j��P�oD�_��_�o� 4��|��JG��e>�H�B)���T�Y�y{�܎��{�ĸ��r͇�K�,���q��/���*���d�����bT�\@fq�5!,���3��;Bd�HM�)�y�=�A��E�YQW��+/�G���%�T1Q�͍|�{��J��A_��͵/��9�.��V��k�@i-,1�g�ۂ��0M�ɏ�$"��4���)��%L��H�F���$�m�R�d~u�VM) �h�jdW�m�T�kvo��*e	��Q=���·6'��r��)�zU�\ߍ��v� �lI�A���9�~r�^�,M���G�>�N���	�g�d��S�?���646�l�'��F	�l@�+�Rn�z����P̓��i�[`����^vL�'ؿCi�"N�ȫ��x���7Ҁ>,4�ԉ��jޕ*}y����M��&�-]����Β�?.�������AB�6w��)n�r-��L_tmfyi�q��y�|d�ƗĉE�ٵZ���L���׻�e���*k/Tv,@�� Ƶr�x�;�ǜ$|�[�B�� �p����:��zJ9KIqn>eV���]��%{��:�F�o$H8*�����W�E�_}������]h���qF������R}�ж��T������#%^�N%�K�vL�ꙍ~,��7C�ܮ�����j���L�p*U᷍���[� �� ����@$}�P�Uo��B-��1[=f��PΞ��V1��6ː����A��Nn��#mHc��($�V��,W=��zKJ�%	��r6�U���a����PU�=?ej@�I�[R}�?��tf�5�jεV�φjT2�y���!�d,1{?����jC�ET���˜:�I��Qw���hp�;bT�s�
Ss�V���H\H�k9�:Ji����M�rOD���{�{��!�=N8�6��/p��Ͼ'bݣ��n���b.A�'��֣�2�5�_k�����5xC-��	��q�.��c��^��2lL�c�3x�-�8�Z<+}0���;/��:�5&�|@����}��S<^�u�`�}	F>*4�ǝT@4�ֶ�0�^����n_�Λ'�����Ga$��GcS
�Iwz@3?lȒ��J���J�Y�n~���P��%�@�"�"�ܐE�u��$�*�+��07.x��.�&�]׭"q�gi�*g�
�(0�0¹�2�b�z?G^ �?��}@��U�o������Y�>O7~��0P�k��X	�_�R�W�*��U��6}�u/��K_<8�|���(~|����m�Y���,oͧ3�ρ��ld�E_�x3X+Ը�6	���o��o`�����C��4Q��Ae�ص�ց��6���R5�@ɭ�Հ�C�/f�`a��׊��1p^�)�1����PJETpH�3d��G3��n-f�	���/��'��jT���h�H�,#��@"-v�A,�W`atv��y+�I�z UO�#�˳j'vw�S��	m;��Ý�F|ߟEɏ��V��3�͐ږjQ	�s!>[���P�@,}E�_	aV�oGqE�2���E�V]4Ѐ����a�$Ǻ�}ND9ڔO�y�7��G�0n�,^h���	7/`�����7�?�X��y(��s
�V��J�@��l��͠b�����Ad^1�{~�qO�}�����qss���O����§�n��"_а�־��*�;/ �e�����U��x�#��&0�-��yC�m�4�q��j/�sE��NG�91�f���l'��3���u|�4}��zzdr��`��N�g�JX��#��d�n^J��wCiF����� ���.��>n�_^~tr�!Sv�L��T�5��zR��u�y�����Ӛ���z�^����D�~�P���j-T�=��J���Ў۰�w��U{\�Cz���Vm�'����Ұg�>ë�Q�#X��3:T
��4��I`���L28(�kk�H�#<	�O��z�����w8w�n'YP�����	��oO���H��[.�Hv3S���t'ղM^�(XB&������A�7C��0�r������'NȜ^6nB땔eO8Hv�&���o�	�Q^������b�v����3��|ob���=��,�|\����r�}%�q��ق/ŀ��$�~X�t�܌.��1~ں.o>σ�V3:����q�Kg�Ω���
�����5QYW� C����M����	A%�o�T5SEeJ�0&���#H{i�#d6��r)���p����6L!?��[����/��ks�^aF�1�.�+�w���K㺎�k���Y'0��m8���[�Kd"���=�hT���������]�Wj���F�p��F1��4ǔKq�}Q��� À�X������ۍځº)рaBx�,Ho�>��S�����؃6�X4�lc�Es������tPP� @`#[�8 #��:����-����1�8� ~��l�bXD��oZ(c�L� ���ᓞռ�1F��Gt`���k*BD+�x�S�?����H+���gSΛs����O󐰅�o@�D��~���;��Hm��m�ے�ˤ'�:�c�j�:�P�FVW�*����죮3����r�%�Z1����faa{�{�vj����y����E;n�h��ܞ��c�p$J�A3�{^vpDNQK3EE��������x�I��m�.��^�R��1�k��.sFJ)�.(73j8�=�u��Um�T�7i�g��<T�?:V�cpaEb1��(F]��$Y��>>����U����$Y��úX�!�����Q�䬚ӕ\trR�	���<�K�D@~Q���.$�cW�xF���7ƠB5*A�����Uȃ��p�����n��i�2�5�6^���v���%�*^�u�t���D�nNcZP�`��h� K�[�m��̙������)o�m7K��PQ�by�D�Q{��s�6��mw~�f���)i?����m�b��#�??~猺�5�5)TR��Wc��#�����Vn��D	љ��.�Y�F�����.�?)� \Ծ����$�Y��h�՟J-~��?®�⣿�m��[�X��\\�~wH��xb@V�R���gK���?�f�^�&YX^�/z�/����1��ٴ̷����J�(7��2����_m�93�|]��.�5{h�!?�7�,�;��ĤC@�Lr�8�Sd�ف�24M*++�ѝAl�<�l6Yr��̷}MD�0�/�)Y5ǃ<����
I[Rr��y2F��9pGb���X��Vw��S��<O��g�}���⹻��;�&.��^�:�"66�����hw}N8a����y���S%�����d;�s���dE*�ǀ�>զ��_�Ua'��k���_����7�֡p9�Oi���g�p0��0�Ø6Ck}`�s��j�C��_�u��A5�R�<C�H����S{��{]gXZx�$�K>��zuK{��|�XlN��"���p�A������L�(�x?�jw0���Pw5"`;�X%�&	l�M^���QFz��{u�Q%�q&�_ۈ:ό�v�쏍į4��B�J�����<_�:\6�$V��Q�|Z�T�J�R�j^d'����'#Օ.e�@amoO����:�N���K����P��]�d��Z�ߺ�F�f�OlJ�pJI�;MC�X;�l���E'�
�sf�J����2��SV���������GY3>� j8��N�B��$8��̇�p��C3�����Ҭ��Եt�A�a[᎝ɍ������W]��]�\'��M��S'�(gE�2�ޟq��l�����^� qA�;��6(⼙pQt�MEN�n#Ib��>�曟� ��i�\��eC�.�膑E�[0� .�2�n'Ik$�=toG[�5�D��`M�r!3۔�$E\j�I�`u�LN�{�{e��fȊu�$�VهY\�,��$�LD�y-(f���ӿ1T���9������O�t��f�Zg��>�	iEx ����[��1����`�зQ���]�o.���CD�m̢� {�2�F4R�8��{��q]��c��w�r�9�ה�\48Sp��򭚭��z�tnl5s1U��L��A�q�
�0�]�y��R�t�	iT<�V��i�C��eP_KΗ ���^�zy��,�J(E�t����6�U�mS�Xj���I�X�.~T�B�l�~.�RZ%�o,���v���5���5����*�bWE�b���:ɾ��#��~��x��P����aL�4[��#�N�ϼ`�����m|���_��0E�0U��ʕ�iL�1�]�r��DP�,0�H~���=��Sғ��l:��!�6XW�k�oJ!�u��ۤ�ΑS����0+�lv1��Z� ��v/,�q�oe��t�����pn�W� ��nC9�Bܗ��b�Xьl ոK����t#D�_&���}���0r��_�J�'��U�����)�
'ʂRH��97������HԀV ������S7Θ�����#�z3Ȃ���1uBe_���ԟ��E3����URy��Y���u�F;����k�z5|b��~��M�gv����2�V<��jثG����yE��\�Nn��D�"Ю������gw��;�G�n�����'t��\gU��/���WM��2����t�h��t9�Ec�ώ��$x?��*{������`YF�����(����Օjk$n�o�kKE]�=�e�gI���T��刦�/���K���~�ĝaHC���G�շ�;Ջ�;#���½��A�rh�il��j�3�"2���|*5�-v��!��ϷV�5���`0+���Ye�y�6���I�-aN�82���@���MYM��;a�.��W�4�&���ՉUz�X�-=48 �xX`Ý�(�n�j)3�G�=&��F�q8v��ڥЋ�v�K����q)�&���0�0K����
�j�Ȃ�]�nNf��i���=K�"�ϲ��2ʞ��1�c��_�+���`8��;�u�=�b)�yr�`�S�47Ta	mX[�͜ڪ	]K.U�o�U[�-����
��uk��,���mB��|Y���)l�2ޢ���73�̆�6��v�gY+�㻔QKD�M:C��gg�+e������z�&9��f+�M�|�]v�XN�Y�
;�����J�GV�h5�Q�`QCL�	�aA��a�e���=x��PoD�y�-dJ�E�[F�&=�4v������]����$�e<U�I6ԕ���j�K;h��LT��}������s!�Ҡ�np��Dc m]��9��T]@�ڏ��^���H7oKR 殿3%��8��.��(
~�� �z�`��R�4��gΜnг�b�D�>S��ԭU�M��r����]Ic>@`-Za(��ة]���y��[S�ͦ� ƯP�=��[~�-Z ���@m��b�>0Xw2"�瓨���R�h�r���1�
�����T�6������bS,��O�&z�&�<h(����?pj�{��n[��6g��$Ȩ��M��)��o�W3R�TܣP^�2�N�����I9K�@��nb��d\������-���|�"���@�;��.ʼH�V���n ��[K�VlAu��%�1#�E[����s�>p�]
��XJ/���Yx4Z�!�	4�#�#y#kZ2Zq�P�|�I��ʓ���c^z��||���#����`!�Uj~�C��,u��N�E��2����J�d�K�"r�I�� |8Kh��>�קN�
��! NydЖ�7��0J�<|�v[��`}$��z� N/�r(<aol	'��`=ف�"��:|�o�q7��=C���|Q4�7�W���	%�朋��F���vu�t�X��T��2T�mn)Y�+WG�5ob��y�_Z�&�}�|�Aa�]������
PA,�7B��t����1�����"���H�`�l�\�(Z�Vi�t�U�5�Idf�p�I�j.��v��v,��,�|rM&˃��+�Y�3*�=��1��j���jX� n�?<@?�VX/4��N�*�X��#���3��Y��F��u]M���>X��s,������l�6���´��G��J.�u�ͱ����f��	_lu�v4������G8�x���Ӫ5�Y�MO��rH��و% �fo>n�:����GU��R5A��O�D	K=�(ly��[���
z~ic�k&�t��N����q���%���He����Um
�y��g��ZT��kj*֍�͸!#�ם6_1��Ǵd����3殱�p$R��^&J�w�-3��~���-����f�Y��n;�,��,)�oM�Lp����3��
�O#���F�d G2�_�y�|��B�� G:�Ѕm�!.q�~ [�8��C}c+:64?���sؕL��ѥ��e7'b�P�,)��l����KO�|Q��,���Gv|�����eE�U4�r�h瑋+
�eN��d�q�6��������X��Т����b�C�~nI��a�d�0��+6^��+�7,������K4$�4��E-7n��v��	O�)z���%L�:s�6ʸ��=[@���|�(7�T�W��"�����N����)cW7���0qEy��K�0�f`}%�s��}1�'4�����;t'DqIgp���񰜏���D񖩽�p��D}�5*8�y��~k��OtŃ���a�(ڧ����)1�Z*X�Ne]��N�OR�No�����j�'�!�ٳjf�H�9�a�S�����'���KbHjb�S�����-��f�.
�Z���ڠs��B��
n�.�A���a>r��ڈ���v���lOg���ٮ�z���T�,��X�E�$XA�������Z�����8�9d�S,ܔ��qbh�l2��������I�O�����a�Ȭ�#JE
��X!tF!���{�Q^���ܢ���(͛��
 �Wépt� �QĻl$�q������~L�'��٢*r�N?�UO�.X�YQ�˰�!i��7�d��� �8��F0�A��F ���X��Wj�W�+.����1�.�8.G�=U�ŧ��ޡ�t�N|G���R�>
�.!>QO�1�������	�5]����	є�a�H�7}��v1P^6�[�f��]��L�j_Ы�:��n?yw�A��v�ڒ�x���[�� XP�`��Q�?���'ٌġ!��`���P�{�B= C��\��w��O.<Z��2s�YI��9"�<�5n�(�C.�L���8�i!�Nv�WĹs���+5揝IWӌ��0Ziþ�(�+D+��5IWI����9��s�Z=��P��!<�#�/g��_���wG�r)���o��Y���{Zh�KL��B�R�*��<��'�b���KRd���U���[�p�Vq���(�`7ԯ��
��?���YP��oa#����a���f=nhIP��D׼[X�JCSL'@�����,�އC�)bC؆�>�ʾ!�O����ƾ�G��B����)3��+��[�:�H�
݄��}�Ue��EL'�$g��>�Xnث:��q- �&��mjS�X�䄿�hg����~.�`s��Ў�g���#J��"?�c��-�d�RQ�NZ�::ˬ��gp8q�BEw��`��������i�1*����KG�BT	<�&WP��u,
�I�/u?�H�k*9��!9�R�Wܠ|RĻ:&v�w&i ���3���>w>2\�G��֥f�$��<7�Z�U�+u�'a0�T���&&ȟ�2i�zŗ���n|v*�ʋ&�l�v�>�8��a� �vA�;ˊ��;��ͯ���?��6�Zc�>K>����w׮�OZ%��l��0ΞıOPg�A�|��}S"S*�ec
"fBV4ķb��Q$v�6;��2�<>��͖#���E�������*EV7��9����F@JJ���@ۈ�/
PW��2��~`D-~`����F�� �=o��g<�<O��c+eQݔ��8z��!��&W*?V:-E��Kه���!��w���!�|5q2��g"Kԛ1a[w��X'�s�t�����h?�k���H���O?�>I��#�f�3/<��z���0_��JJ�����D���8��+Š�CW�j긱��r\� ��Jcy�\p4$�tH@@�����B�{4�㻇�������#m4X���L�=#n����I���U_���Չ4h c3f�w�p!^tމ�����X6=��=$C����o돶���T����$��GNI���N�`p���6P�N����\^*��J��-߆v�J��C�p�� 9˽�x~�n�ܸ��#�[�R�b�C��,�G��<��@;��^kZ5+�"9x_]�zK���z����pִh]�x�|��E���#$B�H�&�9xC/��g%�,Az8��5�-d�����ŋ�ԇ3\^R��,����
xq?xU��af�'���Ӷv�ܧ�2��bwz�59�ٻ����$i�`������r���yv˲��s�X�>�$�h�:J�m��U����`ʫa���u�vn�GV^;��dl�"0���I=f1*�q2�.VTr��(�^���ۥ������Un�[4�'�|6��p]B1%U�r,>:�va,=g��[گ�����i����۲;�Ak�K�v����
<���-�z��6u�J�"�C3TyT:~��Ѐ-n8�o+M���$�ش)�N��L2	�C�P��N~i�;Ĉ�b������/}Fy#y<xZ1ŌMɜ��Y�4��ބ�쪯:8̆U<�~��+@d*o��TJ�vel%	�\pM@�ٍ1�(���3�<�^z�2?��/B��kT�	~\x��~�\u�� ��g@
4y�)Жt6���,�_|��s!��m�Y�p��12ІN:BKyUO��58	k�A�.�3;"�R����I3�Y4-&n������Dw��Zs/r�+6zP	@��	���~��[�f$��� w��~	��� l�ᓋ��z�1���.t�2��I%��`jb�e�f�+v��K�q�����=gc*��DTv������B*�X���d�P��u9��GhJ��`�)��(���3D�<�R1�/����>ĉ�c�W���1ͽ�ɹ�	�����W�DB�3�PM�;l�C�S�N��/�'b �Zd9�Fo�&|�Uj/���E"��߳�����E�z���TE���5�7��/�j��Or�+m�=\�t}Ą)�>���� �� m��W�O��r嚻� I_�� Ǔ���ܘ5цGs	�>"��;�k@ăv3�����1����}t:��Ӛ:~;_D'�LCW�x�̗�_�����c���w!��=N~�(�%��V�+s09\m���.�{Ց���e��&�u*nJN�!���ɯ)*^�r{�����xT���-'tj�iL��p�4R�������8�o'��+\���`��I�?�8k�6��yG�9o������E
�;�n0���\�ՠ��a�_Τ�I{��_4�u	�g,�nQ�l;� _2�P�;�;&'��t�95��3&^վd����{���ǴsU��A�6�n�eC2���x�p��^M=�?!�;��*�u8�"��/�|mh�;"��a&����kՕ<N�]�VWEؒm�d)Gy�I���i��{�$�S[�D�Qf:��Є�|�ցsgm�R�\���jA�C(ʹUR�I�� ��!ߤʍD��h�H	��'8h���B=f��*.l��l����T�(�/��4�{ O�CG«&ZOf���ᶁ��@Cm��Jj��o��=��_z�~
;�J����Q���D��#���7�c�(L��>ʔ�LI-8����^�t�ut��p�����p-rW>�0g�_H�����q{�Ǵ�1���ID[��"�Y�enJ�{��(筗�Y�������-e�)_�-|N���v���,�YWfn�����-T���H����N�j��h׊@TFv"�BcPc��!gR���gF|��@@ ���4$K��I#��-�V�=Ҷ@/��+���otQ���*�x����p^6ɡ���3���-����	lbU��J:��t��鱥� ��!�ӢK~�v�10�����*� &���T��~*g�������:�b9l��''����X^��@Z�[��mS؈y	����_��۔����^n��fT���/���@����?ef��3��s��H��^�H��Ǻi�	Q�xh����G�z��[Y"<���s��qM�<1��-]d9݆ƺݺ�QX\�2Hճ�Щ��.�}���{r$�[���J�X�B+H�������Y�n��w"7/���u��wu�n�Vw!���:(��G ROط�u��A5��d���A���n�v68Q�������$"��0;vi��Eݣ~��T�>!�1�fmL��7�^�G�3Z�Ӣ=l�6E��"��Ƕ�	���"&:^ѿ�i0�K!w���NjY�}�O�eK�"'2%\G�W�ˤg����m6��G���qb?�����`��������f��]aV6�W}�������s߇����r�E�y��B2[d�ٓ�+�LlH�BN=�M���K��"�xr�+�9�E <*i��ֽp�@^�	t��������)m��S�+�}�I���1�M<������;vS���!�U������*�F���N����J� �ci��L�T	���C��v�v�v6&�����;O'2���6E]���~b�f7q*�Ǹ}�&õV���v�|����i*����$>�>nww]�Ŵ�"��U���轏�	Dj�ӳcc�,u��C�I{��(��u.�qtK���Ƨ�p��wK�ɻv�4�M�+��wV��p�]�q�/��p�F�R��l;��ُ�#�X�J�Gb_fE�
�����Աf�3?2�6�(�MDk��Ҥbxfn|r����֭A�TDmlµ���P��Z�~�$��c�+J_�,��i�g�����Z�2��|�6�}�Z���W�@O
� �U&&-�V R�µ���r�E��F闖��q^�!�7&-�>�)��Jł�����,-="^�m��w4)y����e���Ř��N�G`�����W`�KR��.���}%L�\fS����Ln_��&�Q�?�['$�	�xUE�q�o"�L����1�yi�vlr#V�A����.�Rq�f�h1�$���5	I�H=o��BJ��{k�kī-�Ց͍�N���Օ�N����4�	��*�&	��7��^�6���'5�����E~��I^��y��5IM�Ƴ.�`�5���B$Ly1����=��_�����B�)$�S���_4�LЙ�M���~�׏1SO�=<%H~9�SY���6u��� �IϓV~�.�=��{h�0�g���ܷ���|���
����<����@2P9!>\�b�O����DF�@s/6E��V�R�a}�H��
r�^:�<%:��-e���hi���E+WL-�R��s���nI H���rR�����1v�)�ιB��ms�C�8���o�4�/�w|�7�a-�U>�� ��L�`k�P�"�Zm�� b��y�dN������M���&�b}*Sz����WE���	���m�-a�OW�5��
h�20+0z[��Q:�[���+�YħM6��ɦ�����F�4y����t�,�]���S'o�IH�V�3�4�(kc��RA�ݳd�s��}<��H�W����5��$\�>��Y]�-'��a��f��:�u�4������j�y�6���|�X����OjtD�6�>�=�����������L@PG<D��E'�����C�2���F�LP�VwEŦ��#�M)`*�й�J���}��Z���U�_�)�J;uD���uv�a����qY�;����%g�������]��g���$fnU��A�z�Y32�\����l�.��Ӽ�ݻ'���E��W���r�#��tq�h|�s�LD0ꎴ%���_�#��z�-���"u���'�LP�|�˻Tc���wT2v��u 3	)��ʂc�P�Y��)[⩈
^��ؑ���)н�@_Е {�*�ܻ�t�Zd�|O�X�ųI�����+S4q�]�@R�E��Bxu�0e��	�;���@��Y��L�E8��D\C�]`fQ{�S�*u^>'���K�G)��DR������A8\���2Dp��r���0b���&#�`�a�0n�3�a�u]΋&:�����b�`^��wE���]��b��F�ul�����Fk�7�I�~!��u^��i��I�Y���v�W-���hWڏc�%��V��v�޹�	��h�)�רU4TL1�"�Z<?ҩ�-� ۂ,dmi@�M�X����T�	��%�E4--�Q�Ŀ eh3$	�M|<�7��E�oa�۵�Uk�x��~��4�Fm�s�I�$��7\��f��~cNn 䜡r��hR4L��j۹B�ϒm���,q�=�fg���o �.����ح�ue��Ώ�Vv�lA�L�g������&<���ݼ_�o�M)�ㇴ@Q�X�[�V�Ü8�񭶬�7�
A̡���쌑�3)�}1E�E3�r}+JLPR��㞀�R�.t��2�0���
 �Ss��}�d��4U{0�:kH\O}
�p/�4JTqt!�(t[�	�r����*T���^\�%���E��)4���t�l��������>S�5�A�����*`�\�W�+[{�誶�6�cM��(B��s��S��w���9�1z8�D�ŕ�a����K��Om3R�M�}$��..	x��o4����jݐ��*��v?��Yz����O�j�&��;��ԏ�Z:�����\�&a�z�^�ޒt'_!��x�}��pݟ��6OB�CL��׎����B4rH�o�4Y96:Cf|ތ�H
s�i �
XtU%����j�t�l����D�#k�h`��Å�#�"�$�mX�=Z��by>�tv�.ʹ�襀ώ�U�CDǈ��Ϟqx�����[���p���=;��r.0	D]���`� ��7�'c����8����ü�bDEQ�S���b<Z����@��1�s��S��e�ѹ���s�����j��2<+đ�S�b�j^����$� Ⱦ��bX4N��k���A�v�02K���D��GvL�Br|R٬�qwj!lV9b!h`�PhS�@5?�,hL_C�w��y�S�E�2��{G��,T,��*�}�����Z�k�TndZ����Ɨ���z;��"��?�P"��I���Y"����h�C��mS�!��}��f f�9�,Mw8�<����#��y������wa��a\Z�_���2�)Ǝl��f̉?>��A0�P'$t�
�B��lC�R~4X����l���Ww�&h����ͫ�o�L���� �M���t�L[��:,8������"�<������}l��G����1�1O�#�L�+Ts���0�TТ�~q�F�W�k<m�L?Г����(�7Y��t��2ȷ�����%қ�@�]%e��և}��߾)�1�7�g�y�g[�(���p��O9�N��)��@�>��)zH�X�N��,�֟	��¬�%�`ŷ��_��7e�X�(�=��D�~����*�L*yki��q��J��;�f��;1�򒂼.&n�iT\�5{�b_Z��o�e�C�#���.6eI��IS���Olw��������:,D�ٕk�?@ȭ~./w�d�nK9�b[�Ю�������T`���9b{&a2�ew��_!������^�� $0ol�W�/���t���Cً��` ��ot쿯[A�X�s�fB.O��Ѐd�|�(�
�I�)�k��fi�ߵc�_�Cx,�d��<�����_"�O�}B-C�0�� ���&�-����$�:H?ᚍd�W��~w��鋰�n_��Z8J�(z�4�
>?��6���| ��b��h���FI~�w7=�5IWWtݪ�˩a}�%�n��ɟw"�dp0�N��T�%"':w
9����P�n�O� �� ��cS��z3�Z1�9��?�>��;[�Q������d���̵oe"t���V���Ӳ����j%�y[��'Y�;�-�����ޯ��jF�>� �>�6�w/6�B$��A�LQ�HP�h�xs�f(k�F�y\+OE��]C���N��M�;��/�5�|UBI��RuE�	>�g�}����j�Z����3j�����W%8k����zP��w���K`�!h��`ь,]�YR�7����?��^�h�q� �-�.<�?2o�C��jj�_�ݘҭ�(E0��C�_��Ey���`e�t�6����N�{�_��ag�-ֳ7�*LҤ�9��ǵo��e�t�ku£	�K�))���n��"���w���N��#���Q����W����V:�^��$��!f{�i��I�uRr��%���!߾��?%��:���䠭}YJ���'���M�yw����*���M¤V��㉈���GB&d���R�A>����~s�gr��y�)1�z����#5��wm�H�x8�<p��U�P�a�����T"�o�E����1���� �
��Df����9v�#���m��̗`V�*�"g�Up�����ۙ��=uT�щ��7૿�Ϯu���$;6�[7Æ'�\ҽO�- ���zM+�J.B~�(<R��(	�2��r݁�(�Q[R%�ZpG�U�}48�j?��4���p�b8z�tѮ����O<9c�BW,��)�6��d
{����|�	6�frJ_1K��{���D�!��Z� 	Ǚ�DO�` �ɭ}@��,�g�b���K����NA��:���ho�w�]w���]�D��Khb�F�}.e�TN���N�'V��x�E8��r�E��a/�6?�`a��؍N1�j0�q��%Ơ��ɔvH �D;�y��}J��cO��}�3t�����M��,��A!�2�%��;�́\�eDR�pG�2�Z_d>v=�m{��bU�^�$�[#K��"������NZ�$�c����7?Y~��I�k./Q�yh%zp&;����_ �߷��u�����ٔ�2���峓n#\^`�Yj�о�4�M���?���i��L(c�{m�U����r���_���hp�k`M��D٢)��e�9��dX��� Yq'}!�@�`q�S����R�����H�h〓k��Ԟ=-��m#e�ːթ(SpE�$I�.������>�p�Š��G�����|Q�/���,h�}"�x׍��k�?���2�fE�y-OԊ�SI��B�6��Λ^�7J�Q+��$�*˗׌UN8�D�L^p7y����u��Ŷ'_�\[��y&a'�/���%�MI�E|�Ҫ;x��Qi�bD������<����մy����%LXI��+�H�H�:]�]q�0k�\���"��Ť��w�ed��-���� u�蹽�)Y_�h��t�0$h�tQ}��n��7F�4�o�����@G����CQ���"%B��c�qQ��(/��ť��]^�"�_��H�~]	V��]��������0t�"�l�90���9�AA����/��L����6cW�x��X��JO�r�I��&�^b�o^x�z��&G�>����b�s�C?����m������{�t,?Ƕ�ډ�z�Gps���q�D�$��"(c��3O5�upF�� ������ �-�ȥ4�����e�������N���*�J<Ĳ,9tah�W��9|�r��Иt#�R>U~�𱕉�8�HEWkzZj��j�+��Z"ĭ ~[*�p��/�'yǞ�i��Nb�0D�������)��t�{�xF����7�<�6ύ"E����8�m�^�ۅCٺ�H���q�be`�~AO�r	w0�=��r��r�ζeh6���M�aZ&G��A;%O�T��bFk�_�%1�S���W�!y7���d��Ap�u��;�x�rH=SQ�)�1a��=�,ţ�%��eD<Y�CL(n�z4W	�����j4y|�(�EO�:쿗x!�O7������ʃ��okr��7z��<7��'��|!U�F�� �N�X���
r?i�u���5�+Z���p�V����I5Ì5�Q��L� �t�|�Rn4*��A��w�:������y���\� *����/�����il�|n�0���a�����X�H�E�`��%��́O�M<�	蜞@I	��o�Y�7�A��p=hֽ�"��,��U�1����F�����S��(��Ò��E��{#d)�?=uA)�'7]N�b2��X��7,�{�)��e������h�ޓp��-DO���i��ͻ[�K�̻2゗��Yl	�֜.w�!��8�
9=r{�(k����h�΄$�Y쀗Rn�AG�>RZ�.}�INK�@���R6c�,j��B���� �37N�,��Es��<R��-|j���m�5yq��C1諡��R̆�R��l˺�/7�x�y��J{s*2$���&�_�3����5�LT>�lk(�] ��m�ÌU:�@b}�f����ǢD��l�R����(�
�AR��&7�D��O�G��rvyoO^BXm��g�9BC��>�P�02�6�:
Z�~1�؍���2'tR	���HXАu�����1�g�Kh����L����S_��"ߡ|���ْ�9#�h��ˎ�a�S�'����?ӢU=JJ�S~�c���i�#('v���<'���j����K��:��S����6��g��}g��Y	���}z�[��CR�_�k�m�o��!�(������9��3I����-X8����¾k������3�B���m�K�<�� ���J����˝E�H;d-�h�Ph��\S�hQ��7<��F}=|�J�:��긏>0T��IRV�w΋�	T�M�]���v!TcBRN>����f{��M��6�˟��?{�!
|Z��y<�i��~�ˬ�5?�nw�2כ�P7|�[I������ۄ��$=g*hX���"�rim���B�
�7];?�r��)��w�����	a�J��6��mr'X�T^)E�au0�~qL����Skg-t�Ep Ψ�_��C�b(yv���I�,�o����ю�I�:��ͦ� v��ǲ D��j�������ڣ#���vb6��o�hh��?��"0���4|[͏�h�I��q�����JqLe��P_ɤ"5�yë�_A�o�l,0;*B-@L/O�0_Z�Zѩ�ȍ��Cr}\=�4��~-�k�\O1�Iv��N����ے��F١؂�h�JI� �������	��Tg�Z����%؎����y_0�f>�7$;m�x�m%���xY�%2,-�v`8���d�9Nc�� �3���G��'�4TTܤ��NS�狠��-u�� G4���1�&�1��  '��b����p��G�iI�Fk��5����wm:���N>��Y��0~�֣d��v4��� 3G��*a��vĤț�G�#�6\,�s �up"R9�2��U����_`�Q��@����r[��_�FXgt��_�R� �4�d 4V3T5��kty¶ �6$s�6Y�İ�V�Z���?�Nu�C~�C�L�=]�FZu�>o5��-dHb�ltw�U~��ݯ� �Ł<Ȫ�F�x�<��1��mZ�׾v��J=w�K�䋕Lr��ej���KG����$5����o��'L/�s���CS�����m��	z4+u���5��jv܆v��������C���Q�f�3^_ ����Vr�^F�K�b�t����(��	tk�w���%[�V�	�4���o�
\��t�s�kw�����8����D��Y|�TÐN~�i�g����"m<�y.0�;-��XД�"��v1J�uZ�qֺ�ANn�\��	�@yn�=�>�ջ>:(�6�����w:X����PI2�6ߡc�9Ѣ��]�8C��B�k(>�*i��K�*��ֳ�oU�{DA�Lb� ���2�ʚ���&פ^m�����&_ۨ�
��X%<��2z�xo��~�h�{)�[e��5���	)B`��3��f�����(�������kRn�Jg���-a�@둦�D\y'.9�`�,�?�0�_��� �8_�l�c�\C�jiWM��5��'�ʜ�nc6�O�m/5����v1�@A�6`- � �y0f��4��lOEb�S�����۠*��u�T�nc����gL>fDD� xz0�����`s�c�;��!�C�փB�5aZ���J�9	��=N��g��g����-fڅ��L"%����B"K����b�ͼb.nl�qT��)ͭ/Qv݉���>�{�eK�b��
`� IA�)��!x���3��X�_���G���(�?hR����E�q�a����-'}ʫ����^��k�j�j����W�j�. �F��l�츏�^��J�8���K>����_�R?�� ?�c�Hp?=�}����y6Ё�\+���ԳEi�ڝ�n"��96Z��.GD;4h�(�cb(��2�j��#�7Л9���<s�������O�T`�Q�s����C`��k������U��:k6B��$$v�Rѣ��'�o��V�z�{�TrS\:���Js}��\Ƹ�}���z�����J�B�Zo_{�Z޴YQ��2�"��+�p�*�'#D7�p�������1x�4�.���A���>���Nq�Nd�oK��8�a�f�w1﬒��N�'�X�ԗ@��Ƙ��sEXx��?�k�T�W�#|Q#^QNdRzEӝ�0��a"��՜�v]t��{�,�	�bmݍ���E��������+'�L�6�I%�|n��QS�y���W��+/pL��z�T�O�����0PJ㨸M��.��F��n>���
��Jw�Ub
�U��V�-�8�0��W�E.!}�\�="��.�[%����~��)�?������)��V���G���D��j�1`�=��{!�ok)��=,���?����=ǖK[���>@�����$B�Y��ҵ@��ݏ�ǘ��5�ןt�F@`�U�K�+ኮ�C���	���;V/�RU�:���-~���|u( �r,�Uo����@��S�.��RlG��D����P�b7�́�S�"�$s-g֜a��T�* w[`x'�5.+\���I�b�#�|�����|5�Q�\6�;R0;>�^�*AМ�i ���O�P�bZEL�yU�}$��uL$r��LiK��6:��(�̰Xq�],�k��d�:��hJ�m�
j��*�̯^u���AnA�tA嵌��P�cG�A���a���M0�]\L9j����|��lq&9�Й�{NC�Ɵ�g
�4���m��;����lnd�YG>0���Y׏���Dt�j��/$�+�L�9iYk�P�;e�T�a�s��Q���X�����<Q���;��!�t��}�Z��T�e�us*ſ������'"�����8.�Pn����ɜR�fQ���R����ʖ�������O:Y��M�[ʞ���V"!�������w��fL�m�f������M�e��᭼�δ)b1�|���U"�@�?�B��{�����I��0�TD�2�;�X��4�,T=������'��i`�\�����CNiHo��Ϯ��]2��?�K0H���lM�vY��ZQ^�Q5�F�dd=K�_�Z�Z���K"�����n8d�8���W,r�|��ɼD6vb`��]��K�[����ÓP��Ph�����ms,�Ԍ
�QbC��-$��!Æ03��Ҩ�+x4~�v����R�0-I��N/�⣳������~3'���\\e����Rm(�@ur�i���f��(� �aH�����=�	!��� ��L�Z�-�ƤFx�v=q�Cq4^���@q�8��T(��k#�a��畏d>����n���Y%��q ���EMfῂ�e<l�d �Z({ec�B�Gv���1P/H�p�-<.��X,�Z>���~�"Єj���-�#-Pi��+����e�]�A�y�B̍kf��lf�g��eq�d���>{�4\w�K��|X^o��8t���@��XX�o����I��uf���m���jEJ�����4:���S���%�����^�s����e7�k	�pt<��AH�����㪡�JS��]�x��<�Y^e��3����CM�(fȈ�[���o�Pd��:��h�P]T%�D�l㎤
O��P��PZ����.{mG�	�z u��0���SOzw��]��������-��X1����$�r>�8�1Gqk�<���{
����s�K��O�*��h�`��<�<!򘶣�x<1��٧�ę�{	{��$l(W��=iRR��*�QtN�[�(��,j�#�Bh��h��m�F9.���xb�~7�͟�"�2c�ȜUq�@��Zסּ�G����6f��+���]��Y#�&�����uz�:@�B!?)7��`�~L���-	1��]rN�D�@y�yt% ���z��ˀ��u�wQ�7��㒶 ���ڛ1�z_�#ƽ���~�@W a7�c'h	�Ay���&���L�}h�d�뼘Uk�� L*d�,� ���(|�
�_4�	��&�T\�Yυe;��f�: �C��پ�&EUza��+Ϋ�H�k}dU°:���)ԷY���ր"�-d��t{�3�iJ��b���������#���CZ@Vx%Kc��5C۹qv]Z�7,�#�>
�l��OV;��c"�7�u	X)�=!�ۥ�0v�M��8�$���ˬOo�ըB�q|OK�ҝ�1!^7�c����s�] �'�R������Nw'��)����2v���ɮ�ӏ��Ir������?/���̃�y;���0 p�
��	���*�:���kf�������<*\igp�\K�}��y���υ`�F�#	3��f�.-��3��L��:0[(1�
��%&]�B����U2�&;�[��$l`W,��\�/z�����W�tJO��/|Ans�*��M/�M�3'�������u�9�{Ј7����4	���d��(%�r��K�6���^�w��R6���)�o�9z��80
�ñ���?~�O�O|uQ� �zj@�7�Al���x��{�@���Y�[��U��+K"2����:J��bwUX�!G2��~�^�.�:r
L7g�0�uG�RR���.�j���Ʈ�u�&��C��-��pj	Y����C�mK$�O&H��-cY��q��sε�ħW�Q-| Pl�9�$�����N#F��!��e����)B������e=�=�VTe�7}�wԺ�Q��Er��ˎ���0o��<�luZ�o�����~����/�ذ.�)��zr�/�2j��K;�tB0����1�����m�E�4n�[�Irk�1���|���x�F�b�,�:sl����L6���?l��Zg۔��+�MX�,�<��㖐���2Ȟ�,�cX=�da ��Y� n:�4�x��>����Ӂ���$
*4e�4B@�Z�9ݼ����������h6S��Clv�I�o���S���tx;\$�n$�]��Ӄ��D|�9(�	L1����jd�J� Y��%�xW��������"'κ�������
M�����H��fY+9	{��b��Sh�+��0\]��=�����G��[�����1�z9�/sf���8������x�G���A�V0|��{uS�'4��aI'���b�l��������OC�G�C�]$ob���{'s��Q�(����,F�!ű���F�����;�~�H��Wޯ�ĎQ)g�~����O뛦bpVP��\�N��οT+.5o�ٖ��nU[ �a���\p*�� H^L�@�~���'��n�T�w����+n��
���]�
�۳I�J�5s._C�9zn�Ŵw��E�5te��+��LX�*��k>F�*2�T�~�ͩ�R�W�T��K��bQ�Ā����ߒx��?M�|0��Jg͏O���ˢW�>�a�l~��I.�z��ϿX�t��M�_�Z7n؜��	��s&�����W�`�ȗ�)�@�qL2Xh�(�I�4J��+��	�B�����H��G?�<�A����d�*�}π�!+��S�.� eE��u��Ẕ:&9�Y�m*���Z �j�cA�d�`�,�w��A��b���}{1Js���U�^)8���0Ѧ	�,�ɤ����81Ě�e�����������ۑ�?g�`�cnB�,򋙳5hj!� ;��H6�6�%ĉ�*�vNI���AE���<���I3/#��$'�J����(1S�ُͺ7�*,�'�gPIy�'�Ԫl��W>!ډ!m��fk�2��׏bh����� �B� n�,S�[�V���n��p��zs^�5�����o�Т!Z�����E<��Sl��%���<V�(A�8�k��j!)�����ш߹�4j�����5��#�(�\"�?̄�|${�'��Y�|�&��?�o������P�*�|�g��J��ٗ��c�Z�fl�j��g=����!yjÞ	�R��J�0\c�
kٳ$��m��+A+���t-f)���fl�Kx��f&�<���:`��G�A��&Zi���)�]t���<3	t^�lC.�f�����xrM�ԣ��W��Z�O.�=�PQT���o���:A}�Ⱥ=-W�����xˋ��P�	���7���x�K1��zUM�� V��F2�(�d�`ZƎ��I>Ĺ�h���?�?3�&�%��R��K�5h��bY�x�L�x���<�{
e�ʰTf{)�o�s6<dr$P��tLd�"��3^qП�y8'��s�q�A>-C}��[R�?���V"q$)9O������m{o��ʙ�)}c�ȯ>�rJr(��gk�i0/Ð�v}_[��~_�,NH�d� ��*�dNY��8'l��b�r<і���QR�_���l���u���wdlH�N��m�Sfވ�Y�9��>j�����Po�s�DDJ�Z�=��m*#B�0����N=� ċ�ޟ��eT:�G�f<��oR鏮�+l���ƣ-��Pc�ّ�`����O��R/w�u�x�S�	G>q��(m���w����Z�x�RP�0z�ۡn1���W�<PA����=�kBP���7�S�r�7���=p�b+&�x�X��M6"�A_mN�IzT))o�۩"~5��Ȱ��E��F�[�طŴ��Mlj��>� �6| �n 3�	[��$4�Ykk���^�W���M+_��/�S�I̋d���S3���!�.�"t�u��9G;ض����k�y�����_(B(�������lA%Λ;�o�4Gº(X�;���Dǽ���RV���c��*"�C��$YT�Gʳ"J�rf��	��m��ú0�,c�^Wr�/EOXV��#l�Pȍ����� oP]yYk� |Pɱ�����s�_���Jh��wP�̗T�,ik���_bȎkT]��� ��������tɚ����x��,���F��7�����ڳ�	o���|%�]�q�`^�m{]Y-ӳ�%u�?�R3��
���V��T-���.��	b��.�Oi�N�7�F����Ip��<|���	��H�+Ȁ?�߅�Z��b�L�VT�Yl�^�ĝ7�c����S�C�]f�_u��,��`�ǌ���n_����ŵ!wp��T�~X��5����H��f�t�9�B�� �c��n���zN0�Wa)*ɯ�fKP��0������J��.�-5�S�~�@~f�#���;{+�#�r�]�?��/tzbnU��p��j����!1Uv��6`z��fh��5Gs���h��K�����x]���< |����m'6��+�RA; �h���o������^�����"����X3�����O�[	y���5 ڧW?�Ϯ-��!t=e����HfٽH�/4@�܍��L��V4ePɤ*�9<�P��&J���c�~��Z�JKi�ʢ����?�Qǚm:�B�d�5��EV��5�g���h����הp��C���b2������?RP8�����3)�+5�D����n��@��m���$�x��[�^{0�_�Q��:Q-$*��aq�v��s�ݨwG�n�5b��/�g~)H�#x"'�Da��'�S}���O��xQkW�P�cS�Sp�h-�?�y�X�f>I��L�E���#q v�0�Vy�ɋ�i*U
t��&ʠk.���k��t7馩���mb9O�W�\"�#�7���*TR��{YV��\i���a�YϽ@O? ��uGF�X#�th��Jk�����R jy �9�^�T1����*����㿒]p/��lEL��=�F�e������QWo�>쩀�-�z;�2�!�rC�O���v_��f����ʋ��h��n�v����<'� _SLEy�m�y�T�p�_A~}�?��/��RBܩq��+��5�׉��	p��F�]�.O��.�c���I���> ���X�p�:NQ2kJ ���]ȩ*�1��l���*�����cx�T��7�ί��P}���x�݊ʚS���S�*`����,��+@�^�A^$(y������g��O��x�%s���c�(ܕ�� t������E��]�Kk��%VUA[�h6�l�lO�]����B.b\?�Nc.v?$���P�~:�T����'�$��2)�Q��m/q��e�q����fr�M��U3�& �D�(}Ջݼ-4<�/݄����cJuǚR���2ϐ�/��y��u��m�������)��8I�_$�6��H7E篓1���L|6���<�X@���&�&�����Dx�H�y����E4f"sê&%��P�(�>]�!+��8�$.��c�$�g2�Yc�W�p�j�����6���I��v�u�&f gP��r��-��"�$=�C��Ȓ��itA�N�25F�U���;�kWD?a�s�C����ug�D��AR)�Ajw\�O���ɳ}#�v2+�x��n����l]���#��gp�҄Z���3Κp+� �%w<�U������@�l�:���3���_i��P1�D^�5s���fE�6�Ω� =�'���{�[�d�
i�Ťd ����e��?�R��%]�P:��Z�A����N8%�m�q~�ꗌzI[5MDyn�@�`����(�J�I��<���3�3�5�f�yc�M�㻵�sL���m
�B����{����z�j,|M®�E(�D�Y6t@��)q6?�AJ4�V��ٝ1����Y5L�����eF;�l�>���������+��.7�AV�@6�*��A؏�bS[�g�z]K�����r	1x�Ի[�N��rs$ϐ����2���x�'Oc���rAs�����2�.�=�3���I\��>�Ӊ�we�s�߇&�`0h���z����Z'��~��u��=l�̎�.R��H���%��W	��!��:����|�h ���B����c�t���Ű��<W�y����ɼp$���ش ���l6�����|���%�eE��ɯ�^��/*��"~���,
��|���/Vǎ{�̐r���G+�A�u���"��1G^��q�a�6��دڀSad
<M��N�u����?ci�x�X���֧KΦ��H ��Bq���$��1Al��Xg�	m%9h���Rb0_�۬U��{����퓾����9ڶ��`�@۝�eN��c�<�h����F�<���x:�� �����&�t9�ள!J����0��8*�t�^�@�xĠ����G�ϡLɊ��|ʍ��k��A��>M�.�d�Y$	���ӥ�!����:���e����`hd���8fe�fȦ���f�,��0��l��9�~��T����\Ix���Yat�Nt��`��kW���a�F��z�Ʒ�Cƴ�(t�1���,��$��(T =Ԕ{��Ŀ���u�ю;���d�{�1���N��:ciB$�P�Z�x����>gQa���bY���K��oo=��p*@�T`=�3Z끲�^�8�8^C�t����3�^�eA� *O��E�Z�  �;Zg�BҀ�ཁ� �Y�����:T���%81�\�yLU�O�Z��D|z�9��M�"�NT�F=$֝N��kC��~W*�9K�<����F�ItD�8$��6������<�"B����A���F�mm$�6mޡu�Z���25���x�n��k�o�$�\�#G������a�=��sCM�ؔ�THP��X{_-x��#
%�p<o��Qz�����DӮQ ��|@/�Xl	��뉠���<�5��N[]�P�-aW���# ��9d�:�%�����j�P'ˡK,��cu��W��3�|�[}mO5R:�,
/VslX�km޲}r�Xc)��"3�<����-`�ۦXi�va� O���A���P�Q��0CN��ʲv�w�ܓ!�=�~�ZQ#̳��";ՠ�T�n_{c���G��[�]8�x�8
�U��mAV��z��5�9����̃{�"�_�������UP��@������z����@}^����L�6�bg+�������T�C�P�(�]ߵ��a3�$�z���|/nz�M�M�F �� �h>ډ��y˾�gE�8L[��Y��z��_�#��x���c�u"��b�œ��Sj�U�I���9R_��rǨ����`YTo%l����q�s���X�W�3F��t3���[�\h�_�|�*K���"Ν����L�Ƈ�B��W�&�c��5�s��I���G}^}�bQ$r�e٬*����ZX����Ǫ���B~��_H�дL�A���E���:f��)<�vv@��	�k��X؀��a�ٛ?j@|�%�r��;CRJfG��iU�Sp��:��������q����]��a��rn��4E�^����"߭G�^1/Y�"9�Y��QY%b���a������&��l4�Z�7�bʣ�˔��R����/Ӝ;'��»��j�H�X��՗:_4���γ_r���Z�>�R��Ȅf���訩��$-1(c
�݀`���#r�)>7��y<"!���������i��m�)).@RJ��P���ѕ�L��'[z�\8Bn����b.�c�gن	Z�d�A}��y[pM���Ǩ�߭�)��.nQ���be��2���)��� ��yY��j[N�@c2�! )��y^f��[��nba�{Lӌd?�ۦ�|���-��}k����4h��a�9��BCАjh)�g�3����#������ 1�\��[=]�;f�Q`V���N�Ǉ`X�b|X�<�ܺ���N� ^Z�9�6a�<��d�e+�	�0U�eƌg���rc�m�#&�J��N)(eA$B�'�;8�1zɳ���s't����Gw��;Q��Z6��r�?���ܓ����~W�X�G��N�>g����
 b|_��,�Gd�Wu��B�����ɴ�!�,|	@�Y�g��H������;�!�جT��w�1ؿ�����Ϥ3�y�����d�3�W��5�l�e��Z�RG�x�\��9���� �>T���۟H?є�Xo�A'u�Ì�g�C�jZ��;�ѐ�)�dIS��5�A���نD��促�Z���vMZGD�a��BP���	g�.\��!N��t/n/�fP.�Xq�w���_�&��!p�	<�!!}�A
�26��:i��5 ��K�Ao+i2�(���ɘ�
�Ň�g�<�QZ�;����X��\�ߡ�ot�� �!N�L�����W����ć����ȱ���,�CE�qxTA��*e$Z�̠��OQA� 6	e9����!4����o�l�
=j��eF��ݶQ����V]_啜!E67��
qw'T0��a�*�!�����Q���E,ac�;/T�P�fN`�����LbtG�����	m�{k|}I�*5-��`�ֺ����59���k�q[}��{,��'�`��Q΄(H�_���q��u
��A@M���LA�+	��*�г��^���zb�0x��7H�,��Zsnt�6
�;[K�z���@%�C�v��h�7�N^���ˡn�W϶��e�͟iQJG3�ѷ��.��e!e�h�]['.;&�:#���@|�.ҵ�IC�3�a�\���)��h��.aU,(A=>��Q?�n��3>����2C#z^�vщ�/�-�Y���L�R��N}g���4�	o�b�(ˏ]��rI,)۱���W[��?�ߚ�j������TtwaxDIf@J4��){�XS2zs.Y� ��q��#z=
���S�O)@LLh�Ǳ�|��i��`�S�Kz��X�ss|���`���E\�6��˲p\��RҚDr5��^�޲�uwk�:�.�ށ����@\�a�JC�"r�7oo�x�em:�f��f/�^��=�S-��5� '������:ȷ~���¯.�Oehd��lD�݂�VɃm���N(�]t�������L���TG��Z����"#� �w���a�F�㚯��˻�Rw�;��ӭ���S�p��Q��Q�lś����d"��4i�[v���p��zE�>Q=����>���Kp$�e���[�V}GP��d����ͧf�� �u�bT�b�n̛�۽t�ߌ*�f)+���+�ΊD�����({��z9C�I*"�gC���x\��@�(ךU
<5r�3P+�xj�9��S(�_xO��1���f�$]u�����~��Q��|�C�Z+3K��Ř
l��騁�4@��o�W�S���I%
���&1;�3?���h/v#���.�z��l�q��S>I�Boơ�p/:�bD����N_C�[0��%A�^�|�0���8��iypk�8�(�J�v@P3��/����;} �f}J{Gߡ0 .���� xF������/�1bb.r8�jk���Gu��sE�zD�O6�ƿb���;8R��e�ӏ�:�J�^�
颤s�|mt�̗�69��^(a�sn`�uV���M�S��
3�&�� �Zg&e:#�@����]���fV>��н�f���g�D�ұK#�b�O�	
��Z��(B��^��U��8������)ı?U�s0!(I��!"d�VfȆ�D�x���uI;Mv L�w�൝'���xQ���
s��֌vlK�c����co���rI��=�`��g�8C���/���-dt�̡�� �*���#=�\O7�2�}�Z[���n�}ŽW���d�}�6;�cXJXFC�v�q�)\��Bk�P�ϰ)�율����W�,�����v�<�uL��
�����!k�hV�
�8'SN����3d=1�]]ܴ]S1hp��'�d�A��7mDSdQ��ƿS�	8��=�-gR�\�]��wH_�����I)T���h�O��uQ��KdA3�i�f/j��E�����~Hr} ��%�Ƒ_V^X�r��P�����/��r)�2]ƥ�93�u����y\�Ɲ�[W4X���P�o��R�(������e;�D�_������xen��[��s)9K���:�����"� �X(�o�ҥ��}8L��Z(�K�}a�솥u�&�#'.�!@eK�nz�Z��P�Y/��%�4�~%yr�Pg�i@�Ƈkx�)$��^�.|��H��cZ���(����\(�w,��#��z������#�/��d�Y3�d�-m_p�e����>X�y$��~�L;���/���Ho�q��V����� >���N� ���)��� �7l��u��jo��1�)P��^vY]wT�TJ��U�g�~�i�K�_��ȅ=s�����Y2ux���ÆӅ�S]Ⱦm'�BT�<BC��I��"ȑ�����:,nwpu{[`G��d����V�߃{�d��_�h���S��?����D���n������\;u4�R�5�\���s��paOm1�0�*%�`w��lkꄮ!9�9��v L��o!yI��4E�o,U`_Ĉi2�腥7�ل�M�K��AI�����4-�n�)w��O�Ibx/��_-���#�lk��p���|cpCT��u�����%{/��tc�R��G9`��H��x��_C������R����q�HEP���TBVG5�
!8��{-���v,�-�U�Ɔ�.�;�9����0�yN���F��d
�M�E�z��s����<yl`�M�ر�ݙ#r*�$�:�}4+�%ɦ��ƕ������L�&[�	�?W;����v=��t��(�$����e���c�K��-���5��' ����WǱ���6����y��l)�X� �o�Abo���ۿx�ں
��_��|�2߸��Y���G�	��wuq4J�rfn�z��Hᴠ�3pH�ː��h�ԩq�Z��{�(�_���O�����p���;�鹫߹�"&˧�5(�,�C�������R���_�]rg��������C�>0��50�-r#Ik��?-VMLF=k���&�C���U9_6���P�s�6��Ӊw6ŭ́z��K�?�ܫ�+T��mh��lh}�֋��%�1����_����`���r�l��[}K�@����]ȥ�r�Cn���*��,C߬�u���c+�kǒa�@�7��7+��g=��`�ц����8�~O�VOhO�1k���ê�F�gr1�R��Ć�Z��w**Ib߼��;�T�@�<!��g��L�-9F?���!����yk��xk�mԩ�ps˞��]j�!��5�����]/���^P�8�z �oe��ɾ�\`���)C���zo�8��[�֙lbE��(���1�/��I���RTfl�]TKt��Gh�E~� #���]	����>�VL2���s@�I3�~��}P���s�1��-.��` �� kߢ TM�U�G�${M�VN2g��ƳS�s6�@�Or�{�6'BVqt���(�o�1���!~��#JЙm<�y�P�m�빙�����GsϚ��AT؝ָ�iZ${�r����^���n��|�wfj��9Fچ��-�Q�$S�0�Q��$���Ӟ��^f�U�!��A�XbRw�Qd��QG/�
<��kn�We��v�<�0����Ee{���چlQ���Il{C�����p+����כVH�&�=�7hXj�2�h��L��:�����.J�2[m���$L���pZl��(�s�NH�"�wIc^�>	�]�6������q���j���a Ã���acoһ�C:��3���C\ǽ�{��-�q�C����ng�hu���A��a⚅3�:-����XQ5�: �@o~L�x���!�Hy�LZ�ߐ��-�!*,+�Q��Az�hb���:h��&��vU�� �&X�����2^0���|�	��D� �	�Q/o��t�ZqS"��Q��&��jR�W�be�~�@%q�b>����t�U���o�����O�L��R� � �edSk�g,:d/6��=����J�1͏���G�S�a��]5��)�/�Ex���aoD*��2�ʢ͆t>�������C|E�����W�镩�����Y0Xb�<yy��S�z�cY�����z�VM�N���/�28�����6����ye�8�nߘ����|?�T�X#�8���~f�5�_��J�#�L6Jce=y�lDl�0mQYF
���'&�X���
����gn��Q)��f�f���d:I[�� O-�9m�fo��=`���m�� ܸܕrE���>�b%&��;���D�;,O��c�Jt�X{:�`���u�o�Q{�v�iG���d8lZf�;5��}_z� 7ph��ԓIf���X�Q�c�Q��Y3���x�@H�x
�6�ݶ�J��s���؁ȸ�[�q�K�ouFz�P��flː4Hso��y)Ep:v���!ҡg'��u�_����sv��G���M�%q�q����sŹcy�J����ϱ��m���	&W��Y5ï�9�b�� �0u5Jrn&	�íFFBC�;�T�2���ℿ����n֑&OO�f+ƒMzp�b^t�Zd��8tF��k�s4Eϭ<b�H�v�r���=� F���&Yo�4�ܔ�Cp�M��+�v��E�p���"���^�A�!-KjplRp{�,⎞���+z�~_Ǘ�u�FR��D�x��� s�4�E�V�c �;��v�B��6w��Y��N��z�,�*!/���(�ށ���DZ8��^��r�R�4qxF
0�y�)��V:	���f�s�O*�PR���R�����
�@n���3`���=�Lʒ���S��bR����2#v۸�ԁ�P��J!>A`�k �6t���ړ��+����%;n(�ۈ�����@XR�Eu�l6�}Ȕ#, a^��[�^h446[P�y���;Й��BC:2��\�<���E$O����s���~�k�A=7���I획+թJI����:�	��7Mqz�Jz��ơ��d3��]���"n��!��"E�ǆ�6�{��^*��5�G8|P�(��-��l�]#�*]sB�5�2�>����U��.�f��6�I�MM]����1��l��#��X�r�I�i��T1�����g������Gav��@���Ѽ�4�=�[�ϋs2S�Ȍ��_�����g:"M�'�v�h�4ؠ��0�\��4�3Q�K��8CGfXC?{��D��̎����W�� (�����"y����mz#�s�ܙmB���6��c�;ԅ�z@��i��	��d��h3{?��i=M�آ�պԎ/Ѱ��c��7��:7;>�	�.�57�N!�^��l�ۅ:���[L�&KJ��Z�Q*�&���c�u?I��D�I��(��Q$�O����d!bF�R����1�Pz7���gWL<	��I���ƚe�;.5�2֦F0�ƒ�����`��u�`���T�E6ݷ�r<]�;�鰚
ٻ����T�W%�w�N��E�>p��������Kh��G��"<P7����a1h�`ji��S&��ý�y�2�Ϟ㺉�L.�q�Ѷ���y�ſ=x��c��r�F��E�|������� T����E?�a9D�ad���Z��_衣�s���v ���d+��O�d�J�u7����b-ͤ�"v�����e�}$u{�W=;�����QEO�;&|+��q;*� #ŵ(�~�>"#<\I�ˇ&-�J<_i�VPN5�R��w��cUw��-{�mP�&(@mV�@�?��^18���-8d�!���7G�=�RĂ�젤�%>�D|+ҋ{��joG,S��#D��#�yґ����0~�{՛�`X����q	}��M?iV����ѷW�Nɦa���4�S�2�
3���*(�:�S���O>��ak+�"���tNl�a��W�R��e�&#��pS&׆�H�;��T?~��.z��K),���~T%�%^yt$�يzϪ>��w2�S�$���d�U)Y�{�pT�M\?����1 �aya���6Kge��]�Lh���Y}ష2Щ�/��dL��?�^�
2���$�6M�$["n���s�r����U_�06����q;9���э�xA��B�@bI�)*�{��-�}��psL��YAn.�Օ#��"}v��1C�������#�"#b��[FrqR0�EhÁ	3\����M�s���u��A��_E�#�2��3X�C��՝)V�K��fU������%cc��P�M�Va� O�&�0�FQ�ׯ�5��fEu_H��f��MTE�_̵`�v /����uQF"��d�k��$�]�� ���Rw����F��<|ܶ(=B�ByYɹ��v��,ĉ<����i�R ���y�����Bg%)�V�rn�d�εO�>T��N��� W�����Z9$&�H�F5���&1��S#�ӥ`�0�OƆ�ڕp��ڇº�]��2�!Y��GV1�Vt�Q+�9����:���[Ω�hB��p�7�b*u���� v���܄лp���q���aN��zag}��]އ8+I#�+{�ST���P�D]���K�����&���.]<*:Bi¶���R @�x�x`��p�^%���T�d��,N	��eb����<��Y}\�0�P�2r�D̒r
2'��)EO���>Yyj3G���{���	FS�v��&t�'O0�e㩎�[z F[���8e����-vD;Ǫ���1���\K*��k�6�wm-�h��بO<~�Ҝ�P��:��MdM��9Eʙ)�:J�OiCd�6J Eu�cPDd���L�(�%W�l	l8��,�`��-]<�]%M9�Ej�f;��"��ů��,f4l�c�z�����vH6�R{�A����7ھD�;$]�IQ,�rh%�P�ޯ�[��z5Ww�P�����*�2ߩl�D��so�ߔ��{�pf3�G��/\�1�0��뺠M�m$;��mAKF ��k��P��ַ>�ۃ�}��%�r���P 5]uwoY��a�:���0Q`�P��\0�g����sR��gN�M�<lV����2#	�0�>���R�B�^H�_Roh2���Pc�������ю�A�e�  �X��-C�}:�hq�{K���c��������'D�"$�z�X5�R�H�:s89-�O�6d��+k��f�*�{[���k��C�얔���M=�V�ή#!0�߇����{��e�MR?�|��c�m�s5.\`�sz&�A�t���V��5�;�e4��=�tϥ!��V�O���&�lt���IX�`���i;���}�k�{P���ڻ��Q�m�}^�3�0N;Kȍ�C+'��;��]H�c���h�	F���h�	Q�"��HC��������Y�癒jt�豣/)TF-I9W��-IfN&Ŭ� �8=�~0z��C�b�0���Jr�<�oV�w/ȗA����;�����/'���c�W�x.��&@L�p0*ˡf4j^��X=;qD�Y�?�k���Ԛv����F6��J4;�����܏�r� ���g�|�m8��f,5��w�n�Y��	N1�X�^����+!�����q�/[uȼCJ?f����P3Z7��z�)���F��d��)�h�%�F�{�h���>�w:|���U��z?�Şq�?�\�p�kH�xHx:�D��Yx�B�#��3�U�b��6ݑx6�~�8o�mi�i�R�@������S~���\rh�P͕�+6(Á�#r']�����IRZ9~^Ai:=.{ZjL6o�O z��&��]#)�YX}D����E�K��>�,�vz5�z�{u;�>c���4�!��nK?6�yo��{��pȵ�=E^�ux��ċ�_��#4{�d��_V/f�D�Jt�������Pv���?���]�-0�F�x/E֑Kn�����EL�Q�x��8�0��Xm��vZ���as�(���_i6�ja��2d����=�/Q/]�U|9Ww��.˾�N��>t@9��:ՠ�e+���p	�Y%�W���<��k� ��H̕�6w�}g6�yD���� ш�،ͥ��&W߱�x��rWՌD���Z��urʚ֙�F����lP����Y�=b���lO:�&>@�E�6��2����<�_M(��m�~�6�r�d'���c�����o�����=�\�b�=���[p�إj�W)�e:��J��v#I2��'㙼�ͪ���bJ��4�p#!Vf�4ȳ�1�xV��$�͌�?C���0�U�uK��8��o�[�KfbM���H�x�:�2��paa����[�RD�D�E��������d^hM~�#�n<�L�5��l4�Wx�J  ;�<: dZ�?!�hw=��7��Ww�@<�N�^P���s(W���>ڎ�s:��ؙ�U.>W�fh��,��ڙ���1�I�YAQ��kq���x.tL�^�Zn��!6-,�â<���.J��U�rYl����!ۮɎ�/c����t8Y�PK����*�g9IQ��k������}���Q��-K��M�;��ן��m%N��4�b�K���ʐX7{ؾ �H[c��l��!��ʏ#���R|(H�r=��%7-^�q��B�uo�ʊD�I�Ϙ�&����3+���.r2��`�'�e{�́<�t�
t����j*��%ZeKq���ȹ(SkX��c.�b��������* 1�oZ;W�'�L~⥣~[�A�e�
YMD�ڶ��x�/�a���m�GY�����(j�ծ�s̶5����"�4��{h� �&Q�ٌ��C��N�,7K}��m��{�v�F�S4��8���F�.��F��{!������� *�t�=�C砲�ʢ��Mc���u<�24)GN'Ý�>Hd|3B�<�A�j�'�m��M�W����[����4 gm�@��N��mo4]�&U�y4 �B�#��'����j!��
�T����P�~��&K=���~��HIb8܋��Ҩw-��)`�y�*#�wT@G8��%pw��|;6,��h���m�u��*|qd��}� `A.���3�G���R)��t��"H'ٚ��s �5��oių���GM7'~�UUk��q��2	���)����e��"F��@Cy1}�IV��g��,������A������y�v��[X�.����R�b�P��|�Q�R�����%Sі�^�o���ǙPo�di�W+$d���8:ChR�C��{#q�NM��0������I��=�������Q`���ȼV�)*Io�y�Z}3_�_/�k��Y�����'�Go�@�)na�>���w9e���]�ՎSHa���Z�K�����͆eSb�R��^g��Ư�n�]��捻�v|}~)�[�D� �̒�s��v4�}
�V�kh���)��[�E?x�(��s%�(�K�#�E�>��".�8~
���Ԫ��i� 0�!��
�G�(�&���;��C�X�b)l�~k)�/�ЇK_N|.���o�G��~��~�Z;���QJͼY粞P�#i�h(,�<�
���9�Q\��
�ttų y���$>�w��\4�&�F��|�$�^ԡjD�ѩ��$�@���cD�@�
�N��V���?���G��sSH7&:Z��E������o3o5����F*[x����LaG�ʜ>D��9m����jB(4,�M�iH�v��]]�3� L�Ϊ�S��'�T��ʂ�U?�u�Q0�EΉN�0�k���<=~ڸ�lݘ���"Q��'�]���+�"~)P��M�yk���<Din�K �Z���\��i2��;��M��y���JZ��t��o*�o�ng� ^�X�@\�xuG���ASG�8��n(<)����S
�)Ai�'�;RL۞�Q�O��s�ʢ���C�i�% �,~�V}<�hAk8�_}��p�	���0T*�wL7urQ�6
G����Y�kL��`ǚ��6�B���KM'h�%�:)��� �R:�^�a2&�&i�Y�B���Y�W���C�@d��%8F��7�k���,���=�į���͚ī��X��cȰc��A��O�z�g?֬�8Q�^�5%(�g����o '�])ȑ�=�_5�r�o�dV(�y�~P�R�D⼢��<�Q�g��U�*��%Qt�s�9+�1<����,��$�=P�iZW;�J?�ۘð!��O�_�]�ҁ:-�Ιb�N�!��pU1��f����Z�������x{��P)��4�\�D�j�,R2LȒ.����0�J`��Ӕ_��'Ƽ��̐>��B����g��Vj1d(�s�dj5�����Y�2�1�����?K(V[OGc��t���a���1�A��h�rz8�ˏ"1��ؽ��b�0�+�V�I�m�s�GX��>�"V���u�������M���qGr�
Ue�O���{�GW.�z���FDلH�x���c�k$_Ã��}�4U�U�M����EOo�#�-$��卵�}p2�?��~JR8r����.}�-�~�4\zWF��mق'��R��1�>b�U�h��n����G�����jW�aEa��z $���E���6�7��M��P�KE�Wk;&����d�v�����ϻyM������=�U�KQ�ޏx�k�'$�%��b���"��Cf��>Ǯ%��Hu�ͮ��]QqNG�����^c����|��_����г:��$.�VP�ʋ���-d��4���?�bz�n0܆#��RQ�5�^�)���k�m+�^���,�9bB��S`���2n$�֐}6�]8'#��9�],��}�����:��+�}Cy+�w�����u�0Itj1�����"�m���=�2��S��E����������$LUlN���gj>�~��k��-�^�PSe[?*���y�"�,�e��נ:G?rםY�'6҉�x-�uaì�a;���Qq�}���b�hE�5�+/]^C�p������שd[S�Ԡ�<�T��g<����E�p�������&_�Č0s��^�,��Pّ)Y�1*�>���L<�[�������+O����4���%JW#��ya�dl曩�#v���~P�{cq�gT��y*����c�K;�����Y��!����Q��-��I�]:��A��2�+?�B�̨ι���mڽ�%Atq�F�u�Ժ���͛fg	1�R@�ť:��Tv��@/���N~��d�D���?��}��N���(�.>|9�$�5��:P�{����1x���h��H��ޒ O�tC$�A[��ǹ�u��
�&�Y8�ATn�:���$~�;�9o�^͂h��w,Փ6(��=�-�1Z?�=��1_��	�f�8DJk�1����P�0�
_�EgSot�m��z�~�E  ��P4�D�J������Wg4����C�u.	�/}�������=��W͝ �I��q�K��l�8u8���_����n�f�j�Q�a��SS�����'����]n�{���%��v`�������Q/���U��D>oRU���:�7��8o�
��q���ڕ�$��F`Z�ˎ�����#��> ���8i�v�*�P�vL�0�&��U������}9E�z�V����=�u�<xm�Q{����Г�]�]�H���f��섓�F�����ƳYº�OE��*,(,o ��s�"z[�CY��&�4���5��'ʋ�!0��(� Rǌ3sKj�k�w�9~=���|ԡ�-��LA4X�~�pլ1�q��@.3�
��Q�O�ߖe����5���Cgꖏ�G�]w��=¬���1�5"y�m����El�[I�'���4ϠGe��7Z��A>N�uuw��^��O��b��;E	;7#ҁu�cBV��!�|�8 �wqFf��(�Bƈ�Jcָǟ�L5g��&�"c�:f�4�H�6Vn��?�������闓٧/���극�X�Ƚ�#��/9U
��TNO�[��
$B�`_� �����O2�`ⳠZ:@.�i����I�,gZ��8�J��;����<~�����~�r^�]��n(Q��`L�iRGh���-�������,(�&��0�6��N�4 ڠ+
D�C}���P�]8j-�Y�ԉ�O��j�(�ȍ�KD��XH�o�H.C�c?��	w�jl�ǒH�Q�h"�o�h�jM�SId���.!e� A$��х�l���������s,�[�M�x�8�!i��i�dyc��#������]��6�/!�a���UƔD�EQh8#o��͠O(֢��6_h
9���x)~և�|r��Ow#��"�M������WSň�ؒvR�ƕ;��Lo��L?�?<�h3�����+�ӯ:��s��+t�d�����l�'b��7� J�V���~��ad��)�����v\q>�Jª ,]P�M}cm8-�~����X�n�r���azx�Ӟ�����Ƀ�ĤK�j^3�ز��yy��H�*��*��MK�
<R��,,�I���EH�7-}��Ƕks���鮧uM�:h|8po�+�m23^�{4`�c�5Jq�Q�+����3���M��m���j��]j��Թ�s#V�-��]cĂ��1u��&�ym4�VL�M,:�ɖ��A�.��ѹ��;Nj�%G��B�3��9���r�"����qR���4�@�s_�H�P $�Sq��<fE5�����!C�5CF���4+�hi����ĳ��#�v;��B���ҙ/����!�V��+X��ia�ad�N�����N������7�Z]d�>�_�P;7�dK�9T�譱�;A���Ys�ʅn�ܡY,�K�0(�
y�rF�������"V�A��.loca������\P��y2���z�K=LڤiOo�o�Sw��o��녉�}Ծ�L0��<X0��T�ed��`(�o�H�'~�C�t��>�Y
�fY߳�.&K��%��i��B9st��N��78T
pS�����%�8u$4��)�n���6)��k�u��<�@��I��·2 �|����̥	Ǖ*�>�?Ǽ�r� h��������)�XA�]ҁ���mݖC�V:�E��v��m�!UA<��ƕ2��7�:ո�j��1ゥ��Xr`�E�Z�2����;+�B ۏ�{��I9Ҹ��P���b��ϸC�e$p͇�����?"wE�;�*��B�!�1.Q������3������dPޮ7*�V#Rk�R^�n�}H��#n����޽��G� ����G�P����z�WPP�F��!�RS\�V�����]��$�4�EF`�Y�U���z�7�~��t�en��ǳ�pQ;/�E���e�t�͛�Ij�J�˴՚�׭7��I�&�F	���R��*��m9���$U��+c�c�.���&q���L��bE�n�E���]<%�J��ǧ��zL���p��W���"�� %�^�r�JT��+n_����?&Hs8Ij��R�.ڿ�~�X���82��Q&rJ͗)y�-G�;+Y�п�X{Z���)�~6*A�*�p|>�x-���.�u&��0*��󐺢s۟�5z��i�q���t<63���vn�G,L�7�B8UZr+�����˛%���Q17saג�
����5�q�`��J��zʰk��a����.xV-���e�9TA;��W$i@j���U�&��P-0�rm;����C���r����=)�L�8dt��-guvdE����@�&_9x*E(8�b�>��袽h����#�V+�ﯵI�Q��R��P�x|�0;���D���SPr���0'D�u0�����N�9��OG�<و�� �2��Uu�_><%�UR{������� �xl��H����Yqs/5փj+�爿����F%�e��c㪢ϬW��L��W�i3��q������
�����JO���Vh�	�I��8J�5w��_���Z�p���m��R05��C{Lsp�Y;�C�&yq�7\E7�נ�c�&I�bK�!ԦA�m�0�'�����NT4�F�Q�PM%v��ȁ�(�l�ʍ��Xo�;b�tQ�L} ��_.vc����a�4w^go�`պ��4��oϹ�p˷&<� �z�z#��I8���K��{8R�:���T*b�,*pnG=6�wh��=���?�D�y��}���[$Q�E��3�PO�w*"�f󄀟�Е�4}g�Rj�6�fD�Ň��V޿L�)�c�(���"[��NՁz����W�C�=XN��G�)"Hv>{�>S`���9���0��^�q���Y��Ǻ��ѿ���������L�qiY�J���+X��>��wๅ��+�-�`��E��DQq�v���i��{��Ǝse1sRb�Z���|Lc��D�?i-� Y��ur'S{�])��r%*�a�����4��p��"�frv�n�Bem�pu!6�}5�zOө'��"E6�|KA
���N�xf����-��͓��B�!�ds������Y#?�m�����1b���&?!�I�	���9����/ݳ7��0�_�.��R3�h�˿SE�r01ms�1I���>�q����� ��`��)|�}8�@����T��!<�?�Z]Vf� ���Z�a�?����޳��3K���YFEp���V��d�[p�Q��SqZR�������ΠPh��v�y�n�-�n�LC�MY&>�.N<���Ē�g���W��6��ㅹ	�N��U�C_��M��n�F���gG��@�*�t�Ā�"ƳM
{���|{�g���)��(ȗL�V$���>�٥���xʡT�dTZ��N�{��1o"0���X�b�>����H4�x�Z����P��J�_���K�0�^\�`�>�����?��Z�s�sy��Gz쇁ԕ�ט�U��"�W�)ҩ��;d�ۧ%/l���A6�k�DXI/D�	�n�1m���N섄���B%���;�M� #��5a�ʢ$���΂ۏ�p��;oo�9_r`Y�>r�4�1�6�23�<I��y'�����R.��p�*-&�ږ��8b���l4�@m�a<��Z+�������9>K� ���G����۝&�C��1e���e����7+C
SWr
�ꢰ� w�;#B��`m��ii�r����
9�f����;k���Y�t��(Z,��g��wT�1B-�,C�{3y?��LI������<.e�N�0�G��R�b��N�#�R֥Wz��E=�HS/��?� v��F�����|T8	N�تlk�J��c��6�4���[?�4�y�)�͝�z�2� ���x1-�3u����a�D���z�p����������9k�V�GQ4�&fۼ=��ul�[Fr%$Ή��z���E��B,�(4|o;`����~���#� VL�-f�܌ԭ�E4=��Y�i�M������eb����t<[�A ui�9�9�b3a![�VI���ft�[�͙��ζQv�J�MI��&e���)J�v�����͛��N��*���|vw�K�
��89yq�ҟ^g��YB�9P�'Ȑ�f�A�9�z�W(
�����%����.�V�\Q�ʤ�n�:�A�����cD��p#��c`Wщ���l3� �FR�E3�۬ndk�OH��6=U�)6cX����i ���T�[�}X�j\�,q����w��`$�H�
�7]\#r����W����߄lҭe�w���|3�w�>g�_8�/w���f���p�!HB �9@:�"f�l)�6��I��m��R9I�J��З�`�"��D�/�����oP�}�۠Z�!Y]|�����".WW8��}����Q�
�����S1��	�~'4�r�/厌��e'���� �v1牬�қ�Pf���aZ�Ūx�=l�p/��R����D��kÝ��2� �wN�m��)9T�Vk�\��kS"�����5�@f`M�����pp! �Zz��
�4��w�I}�?��]����<�%�P����_�Xܡ�/6y?�ֱ�-��0R�s���moU0��g��̃ϑ��C&����Y:��K1F+��גXr�Թ���'b��r+˅�_� 	����\���틞Ν�+	���5Ǥ�E�/�{TO1��;�E�M���M0���sU�Mֿ��6Ӽ���ͪ�|Ktg�K��5���%��}x-�j��I��@f(�O��-0�q�3\�&�UBgPv2,���:Q�ްi��\ލ�=�,Ъ)��Ès�л:cKH$�@w��U@����S��.�8z��I0ũ�۝ܣ6��Z<�a'ݻN^�jVm���`���<��,ad^|�&�I���*���i�2dp#/8���}*��R�:{�^ؒ��+���~�P��Sk�����÷�P j:]@!U)M1����ç�5o�t����#T'�2ȭ����m7����v�s�n�<�8poRI3�V0*�!�T�������]��s��J���:�>j�W�m+}��/\2�;�Q�� 6ő;�7��#��eߌ^3\��
C�esn�E>�ܱQ�k�(A��>��/fD:M-���"B*��@͐(�4$�o�X�~X�]N�Ë���N�d��l��BŠ��@r����W�����K^g���ChT�5Cm������=���W���zi�ry@�Rku�ZXQ�HAQ���s�>WV�����o��L��;Z	O;�e��'��Un|�Ç�4cϏ����e2T��J�(�M���J���:e�Y�Y�� �Y�D9���o��ٿ�:� 2d@Ṁ�9�;���Y�o�����;>Q��p��\[����'�2Θ��:�y�%H�s���2�s�cM���wt���l����Z��_fi)�ohi�a��z-6��og]��M'���7Kl�T���ju�2:�D+���BT"� �Ƭ=W�i����ͨ�*��u�ڕ�Nҍ@�P��+]�������G@�X��qb����"�J�h&�n2g^!�>��) �v��A��L�	W��kv׼w�IZs6A���T?Y.���*`�S�K��9m�(=�EI��4~�u�_u,������p�����a�^�ď�D,�0�82I�W�{�ċ��q6�!\<�b��*�J��s 1L���U�Q˩�ƾ*��6��f�Kb��t�i�V���r�Dg�P4�|�~���B��e����W��
�q��y	�����͘�͜8�ڔ5���sH���)��(w�r G��0��,.qD g
�ךc]*��!��Ez��r
t*&{;g�3��7��Ğ��^PS��_2}[mC��a�)��I<U�Vn���5�f����q��dy�_��>��/��8�+]<+�u���%����m $	�]9"�Qߍğ�:�:E�^P=|���+��<�##�w�J���xꆠ0�����8X��Ap'�F������b>��(_Ĺ	�(7��dT���.tE"��Wyl��%��</d����Є��t,���@
�)D~+;�NEK�"zGGq�hFh��I�l�	��^Fi�4Q��u�7
�.rQ��H��¹f��b##��� V��L��t��6Ґ��-�=m�lӔ�� yS50���p��Z'-��I&�=EL5�2�D��6v�Umﯹ�f��"�&��{��u@�?�k8����`H"�]�$%�cp�j2%%c�-�o���Ǯ��˖��4u�&�6�"^Kw�w	��w(a�%���:uG+��������Ϛ��nߚ����c��y�ʩ�������:edwg_P?�LtU���<j�&jOȳ�iNC}E�,N����uN��i�ք����c��110��]ӣ��Tf+��'�xO�P�<���)�gˊ�pVF�7�i1�����',��#
̓h�+a�i��ٗո�Z����ȱr��+k�N]&���A�a�-<=��ƝF��YVx���E�nuȳ�%\�L��Qs�v�WO
���~9g*�ƻ)u�z�*��k�o��O�S	^�`���GE��YP��3T�wEs/�&���j��v�4�5�޵����k)Җ��r$G�j�ݡ⟘��ClE�N5ao]l�~����cr��l������ʰ�'���x�73�Q/4��?��]��vH߽�zt����k����%T��L�_�\��l,?�t((W��{��kp��̀5�vH�W3',�s�>(�韂������l^���Ҥ��k��ݥ�.���ɯL=�4�O���E�Ofk���vߡaɧ�ē:)vZ�E�:�#̺�����UCV��j��Q0��h��6?/w����M�I��jK� �CF�îC�w��8e<[����C�g<�$�#M��Tw4�);�2�\0r�lOʤ!�C7��8��{��L��׺V��Ք�:�:X�J@a� $#.Dm��q|LH�*���9��㊖n��=�s���3�w���w��R{p�.��Z��o��֥��Q�K�j��J�e��}��au��|Z�=����0�,�RՍ�L�׋oN ��F�|�K;f���<(P�␂H�z����&��Gb�t��Y<u��	������j��t�$����lo��l(��Zy���LC�K!���yמn��%M��wq�f[|K�(�e���[��u�p�6w�aӧ��?��9�?��F2;�}�s|Hy��W�h�����l�_=�W9�|92�d��
W;�IB/���Y{�U��<rM�0!��g(K��?c�����y�31��I�Q�Ӆ���
�X��ro�U�0~g�W��T�-l|��]�C����1$�@�@��=2�i3mܜ���Z��Ϧ%��ߛ���	�r��Di`w�/f|�t���$~&�*e�/*�*�+.ɖ
`���氡����.��I��BM�y�Y��뮛y�T!c2� i�T|�@��~�X��p$ Ʉ"��}�1��e����s� C��p-#i�~.j��Gqd�����V�{w����J��(��V]�>,�B_����0jo� |,��,K�㚊%'NВ@�W���Y�	�H��/w�>"-�s5ZRI��q���"�C�x��ɩG|w��<H���˟QN�+#(����o�����P�Yv�g�@.ԃv
����H� ���e���d�2�	m�4U�%�$�δӥ"9�D��Q�aΕ1�pZ���1ro���XkD(l*���{�����)�<z�hib��"�9d�XRLԏ��gp[ j��Pt�*> x�MdN�t�N�.&�� [�5TU�d�Քl�(��R�'�Q��m��zє��FO�UM���qƹ�B9�Q��uT��$?ͻ�9kq��&���/5����P`�H��m�&�?[���A�7��S�n=�7C�7����wd��_����-��x�#��ر��SRs/[i��$�1��^tvH�6wqW�b����Ј�D��Zl���X �L�3s:�f���С�����oFF����qZ�A�k�6[˽v�� Ttts�l1�؎.�b����x?�H̺D��1_��o�\�H��KDH�*�Фfv ���A/H=��R�3�[�؏����e/�`�Xq"� �0�c�Oi����*���.%26�吙�3
=�_��n���P�G��*E�V?--�.�Ĝr1�'��C��e�/��x<�,�a�16�#��u�_2Z<��D����O��Y~�`d���4Q����@��t����V#Бƛ.cB|�[1fA����9��+�.5�-��%����Sa�ec}3���i7�h+,�EM��'Rm�ѱ��ᒗ��a�^9\�`B
����Df�z�������gJ�t��z @�iGvֶ<Q� m�1ڜkRؾ֤u�f.� 	��#?���N�L�����yq����i��_*��"HY��^=L�>���Xxv�>��^ze���"�(���异���?op�����2FE�ڔ�<XC�.T79(�v�!&���^r]�\�E��C#ڢaS�.i����̏���u�4`3��F��*()��S�W��Gdz
̯�;f�K����|k�f�5��,M��M���P���T�Wց`��C�w��`�t'��?0�r���mNV���iwSMBJWb���8+Mގ�p+��Դ1겶�J@�ܬ��s<[��`w;8�Ȉ�ѐ�|xQ蹠5ъ���7��A�w×�B�W�ެ�}[�bb^��G�N��~�5���*l>Z�q��ߥ�0/*w电����`���sEW܏��T�3o�|>0�c�l���}`J�i}�`��xI��C���PCL�jH+��d$�3�6+}UA.09���LBk�-�z2��t�����-��k�x�~V&p(��Ѷ--� ����,O�	�jX�/M]M�_�k����?�Ν	����SMJr��6��Q���s��~Dw(��g|��('�軽H XQ�	�,��.����.������*=;{��{Y�	�4҇88u�c�Kjq�mvA�a�$aO�5<x9�a����n:_�+dnus�H{��7FD�6D�~
`��ۨg�6��'��*�xR��h�7�{�A�ا�5/��Q��ۺ��+���P�}�/Y��4 ��L����_irXJٚH���^( ��`�վ�N�M1�SD����q�����5r�J��{~ܖA��6EMΗ/��������e�D�����a��zԭNV����W�K|�p4{?r���P�t^�yedb3�~�]E{<�{ %�b��������v�t�&��b?��;R1��V}�4��H��ы
��?��Cϻ����_�>Fd��*!β�f��9c��o$
ҼkV��9�z���l���Ic'H���;�)�+hBt��uS��v��Bm���W����K�5���V,�1bU�q����@�<i���.���<��Ҭ�r�k��`N�i���g�0!gt�7,���Xcp�Gh����%2����ME!��z�x���$l\�����M���8z#�������*����ٷ�m�9�=Wb,��N�H'���bEa�װ�r��3_��ymJ�Z��29�!��x|�a̐�qq�P���ӕ^SD�C�>�ʷ܂4�R [3�{ޱf�=߁�!֓�}{���[VڐoߜװH�|7l�FT�D��'ٸ������6`��c/s�g��b�:f=px�->n}�u�"*�w;sD�>�'GF��K^F�~2�t		B�6��̸�F?P�`�I@�6�Hk�DQ@ݜ���ӻg�V�9gr�8T�m9���36�o�ڜ�D�у��7v¶��"�Z�2L�O4+����A?v��B�ebo��J��
�j��;��$,�.)!�]���ƨ���7�^�������e�����й���1��֠��]x�sSt�~V��a|zv ��n�b����E�̞���f���m���K.��{ݭ8P�8��7�q��>�A�L�����uh&&���@R{qZ��ahD���u�~���H䃽F��+��Z��Å�:�&��D�eX��uL�����9�G�A��?h���P,/jҀ�	��F(�9oRM�8bf�t�+#L<ki�Y�V�Bm�^�E��������O.�{c fO�X"I�M���>K�@R��7��%�;�b �]$~��4Wy9��q�^}�*�Pfmm)F��;+]���Aд��Ü+K�D5�A�lXW�߅�ʣ@����vn�ՒGR���z剐�V��<2�S�)�\�<���ӣ]��zGt�I>N�L�1��Y���<��5.j��镸'����Μ|�8-H��>*>�\ɔ����N�F8=e@мGl����T#�Y�0W=5�ζM$5��ʀ�Ì�:y$�7�_n���Щc5��7S ����UOWr�;��P���TS�!�B�{Ap`��L�w����/�`�ۑ��~f�Cj��q˹��/x�S�B�fɺ/&f,��Ӯ=8���	�	��X`~�<f��|��7���(]p{��'恂i�A��؋b�E�"S&���/y"]#t�9��ѭʜ9yG_O��t���t�9ݝӣ�:�d>�2	�n��ė�n��p�W?U��6?�[@f���~rh�dI�ݽ��h�R=$)�V|�� �Ɛ
�G7A��;�K���u�:�7L��sx��ӗ�S��AJ�q6��;�1�bx��,++{��Z�<�ER�N�y��*i߄h=A���d;i�^�㖄�3z>{��w�(niO�]8�+"I���.�h����Nj���Zdo5�����}�|c�f�((�����ղ����&�Y]�fsO?��N6���@�՗|p�)������C�L�L��/�������=������j`���)˚�7�M!�v]��>:��q7Dlր�Q�g�z�M�*V&{ Ai��ѵ��.XX��[�9+����Z9����G����I�U��O�F�}�Sl|.�{�q����X���l$��0�� e�s J,����M5`����8��y�e����
=8g�0m͞>�b��*5��Jh��#����Y�����φ"�ҥ�垩o8��k���I�>�{�����8�1f�P�h�!wm����0��s��t��`�Ib�#�/���]�M�U�K|�-�(�_�R�����6�3��q')?�̶���w4�`gx�Ā�B�vF�nў���~�`�st�@��d�~�JQ�$��@�ݻ���t��D|:�)ى�v'�j<J/�꩷B3>|<:e�"E�[�ճ��~B⚦7̀%���D{�9�v* 4?�^�ƣQ��_
auo]��P���|&��m_ ��l����f�\<r;�t=�(���{r������	_���}�kꔇN���"���)�&5�e���~ԭ���1�����2����lk��V��K��d_�}�<��O%>$�R�4Y�#=�l_�]��������iz�+tK�$}\���K�6|��V�-]�幓���6�p�~T�R��1߬$_��и�_U\���d����,6w�3�V��_g��#���w�-ori�*��6�L�GyPo�1�05w�B�̗���X{��r���X:^.���{F ��D*�ĬY�^�2�c
d�f��r��z�v��Όy�����VlT�z��}�|Y�z��9�%4i�P����y�(��vṫ��W�r�V�!��f�;�0i�L?�z�V�a Ŕ%����a�(͓�q����AN���: 2퉁�?���a�"�u�9���2����d�m5<ϊ��s��
V,�hF��[�X�H%��"9�v�l��+�$R����>ޜ�	d��8~���F}I�G�m�ݭ�M�F�i׀{�}�\'�,}��$���[S`JH��dA�J���� c�S+._��H���g2q�8����K��z\ؿ!U_Ϯ�2�:b���P����z0��������!Z���L�IJt�������IjFftd �}����ť2)q?�ɬf0��*j�o�ZWm��#�W���NY�%<e*�:M�����������,��}��m������:>I���ș��bT�|�՞�'�-gQf�q�Y�X��/����:�G���~_hd�!�1F͈���j,���0���)�ي��w}�!�ܜ���n��X\׋�߬�[˘�v>]З�u����K��0�DX��au*)z�U�̉�����ӈS	C��Y��&�l��g/��Ԇ���Ysm�0)���O�����̀��F���~�����Uu�T�C�z8��'�!ƹ�V\��b��A0�{����Ph��)U<��eCCJ�4"C�
�nŘX.'����gB#d�T���mDO�4�b �R�5(b�N�<>�ߏǙZ�!nQ�O~ �C����������b���8��2l�O>��NȲQg\6�$�h�;�hg_�q��Oe�6�2V�����C���Uޕ=@����G3���=�,Q�;l��FZ���d� Z���y�=�=����s�����1<�:������*�A+�H�+��-����|:\O��/�>U�F��GU.]��۵�-)wK�!���`�ew��g
���0�nOG�����c�#u��{O�-�K*Q�� � ���R�x]�Qսp�8�aHk�{�����-�/S��Ceź�풯�W�4ա�~Xi�*�D�b�����Ppt�)��Ƴ�r�E����vc��(6��A���0��۰غc-�>y������/��%�<NK<�����ț.��
UP��K�{�V���-!{;�)�S �r�4���[q-�Y(%�&�I����r/LYVi���L��D�@�AB��yu��t?4��j���d��7�<�1X�%�������|�\�)�u���N`��M\��D�G�����C`e��aW�w�H�a.7���_�j��K����5&=���L���ڇe~�����r�U�J�< @�slI��*c��~���ͱ����f��ـ=A�~�S��id��)f�r��w��+pt¸���.\cg�#|۩��2�!�NJp�3��� ��Z�I.�Y`Z�H-w!�T����� ��RYX�7�	Zֻ�*�a�V��=�N/����B�}~,u�K��;{�T@����r�*<m�I�hfְ�n�隤qPj�8b�m򑌖��&uopg���g�Y�y\��öV�u�O:B'Oax@��ܼb[��إ�#����d��C��	J�첬p�D�h���ͮre&�T0���q~I){V@9P#��
�!��`�o��﯍��~�x��w�b6�8��ఉ�[�@Hx��)κ����!3��T%��Ng44m��n=W�ވP;�w��^�z�o��ڵ��N�_���p�]�xq��w�!�ڭ5�C�h�C�%/�juяMrN��Y����k�SА-�R>��nfU�x�Q��������Zv���&d�\��Yo�2l��fm�e&d����\��K~������g@��t{׃�̠� oӰ����߫�a��A	�y}.':����*�2Ca�,O�USaG�꜏qLܖ��8Š!�V���Fs�lp���w%�K�>��,a��;�x#�o�C��\�����-������9�P� ־X��=�.��3b��c-G��Ҽ2�m�L�{��+��C�eV�n�����n�s�H��7�d<-)K�z�
@�)i�T4Z�S�>Ni���D�U'�|��|<ht4|�м��������Б*���{&�홳^�90���G�ɵ��^�l��{v���w霷1�S�^�k���"��G	kTl(�����I\%/��q�BK���������"�I޲[�o�U���	�K���4�un��#�1�Ե��2fߌ;b��G�."��#���ʪN��X14/3AE�;����:Z�,�$$�̍�Β�2M� ��͕8�����������_S7s�{O��L�S'�ʥcW���d�
��,���rX-?PVB�������M�G�T�
,{�q��ٖj���,�.a����o����~�*�|jb���e�	'<caߥw,�i�"��t�v��S������������ʍ)��Nt���Cob�JX�R�bA��`0�m�@ku���}�J�Y��zV�l��
ʳ�ꭀ�=b�g�3��U��l��%�݃�ԫ焈��0���u!����i��K��Y�J:T!�0�G�1r��D�q+��_c�8?G�f��鏎6��Rs��Q�����?iH1>�6Pǣ~���bU��蟿O�X6Η7J1����������e|_5��>6��γ.�.�	�M����Enemـ+���|�k�QWE��0���,��� ��Tٟ��h���si
y��Է5�$$QO���!
��tRb�d9"ܟ�`�NQ���%D-��u�I�w[=���w�/��pJ_���6�������h2)I��:�e"��V�)�aJp+vυ	j6z��m���S�f���<�	*`o�����x��h�B���V��e������#���?�4�O5	2b��#���ޟ-8��Y"ZҪ�z]�%;�'X��[LṚ���1.�]�2d�t�.�<�pRQҭ�m$�8Szj1x��Ma����4�+�K-+? -�5'��h���@u�]�dNs
'��~��2�*r�=���m%;%�Ce��R�>���<0!^)����cwQ�;�����UY�YRW]��JU�+���&��+'x�gF�Ϟ�4�RWə�A ,���(E`E��̒]�������u'.�B���X��D�M���]����	�ٜ��X9�K[&�i�p���ޮ&q�aZ�&H�o���_����q�kC-ؗ�c�:�W+�E��^tmf1%�Ф�f����`�q���:�K����bN����@ՊR�f^�ޔ9T���j�s��q��{ g��� G%��:��g�+�>�bؖ���m�pѴ�d�� �&�u��1f�"�z$���#�+ծ����f03/&q��Mُ� Rf����I&�S���s�Y��5z��D�bd����J5"��0�� ��URǚ�x_M'���w�2Ԏ��(��f3�������)�Z��(hu��#��+�)_�6�����Zxҥ�7��̿�U ��э0]@��J@���a���e��}��96뜑5�~����'KV���񂶳�Gx�%��e�_y���I&,�`�w�Ő��]��jzvD<JU֑���/&�ly���r�#���'�����un0����F��;�Z��a.��n�&Ɋ�[��[k�,����X�	��l���" ���K����pAk�/�r���M�#a�L�٪��0&쮨Ќ5=˲OG�}1�x۔�h�����y�ai���3����"劻�%r]d�@;z��]˺�[��%�U�T�Oy�C�B��Ud�>�$�6�6�ʒ�������QM��?-�������}�q���~S^r���<�>
�s&=��аY��;9����8+�0�)t��+�h2�1]������T�K����i4O���^�T*,�'h&1Cmph���]+�M��o�F�;����ej�����C��_~LÛy�S��oqB=1y�Fy�9���ݣ��w�V����h�1�<$��j���[��T;q�O�k
	��r/+.���'�5���g�uz�Aq:zc� A�c�uW�tQx��@��8��O�ޡ!��Yye�� ��~&6�j�?�1��_��X�W���R��+��]x 	M
��҆�W�ua��2���.������X$��X��vx��*&}���LV�IT#��$Ƿ�F �}�M��Y�X�%\|�n(��!3�5�Z��f=������q�y�e�F
};�h���p�(�9�2E�^GF��߱zn-M��~&� �e-�O�L
Se+Ɩ���:�︩��RLzJ[|�(�'�<�3�]�XoB�寥����`�e����A��!Y��&e-c'zP� �o��y�f�)S��3��F�<5uq�/k�����e��0r�?����9E�
�p2B���K2"�&��B*Ü6K���ha�����bV��&�:����9����Y�s�T{�ekQ��祒�8����ەϟ-���.6Dy)�%�C3��@��7e�,�Gv0��.1�/�xfL�����OI�X	o��q[!)������B~c����F�*�$5��Fb�[��"��lt:�F-��zL�:�VүO��G�d��?e��d�3�0�4v~:�n��Fu��˩�%�%��t#Ҧ5�N[^4+m��1�>~�6�,Ϣ��'�36Zi&{�
�_eVZȋ�ۨ<_B�aU�ӷ�0Oʌ`�;�vC�ӊ`t���o�����y��R�M��0�\�!�9s��4��W �������%��^��2�bRn	�[��G��kk��g-I�e�$5NS������(���6V��a���)[��K���0(�Ƅ�x�ƈ�Mu�V�z�0[�L��kKZ��U�0�f��	��8�k��eByc��D�ˆc_�O��|B����V�Hg�|������S`�x4Q��88銬)Go���l	���i� ���	s�o�"����쒬Ф�s���rٙTt�t�:)lb�n��<v;	���m\q�{��۹���!�kDs�1xFZB����(�D[�A"���w%cM�Z Æ��$,�,�������"�x�ƶ�����\�d���|����	�D�Q.�����V�U���F3�2�?Q�K��"4��$ЇĄ�&e�i|db�'�^����;�P�~��ϱxZ����М嶦�=BL޹��Dg���b���tk5`��u�^�A>֬���}:�� �4))!����cS�E\w�[�sL��q�^�V�SCc��ۄ	+3�\��Zn?��%��R��̟H�=\L�\�rZ��,<X�<�����:V
3#���mO6�%��5�����.fG
�vѥ$n��E�B���}'[�۝P�� }C����@�G����Y6ԥX��f
8�m0[�S��C�@�?]��8����kb&�R;%|X��7p�����I��ϸ�t�V�0ކ����Y�l��p x^��!��]kC�s�΅-9����gb��Рj5�M3���UǨ�7cR��lw �-Gʓ����:��Ͽ����w-@��(�kG�@D�3PL]�&�d��	%aL����C���S�)��D@�p3��@�O����Щ����0���0*�J3��A�|;�$a���{
#�`v�0��ѻ�#��u��~A��>�O[��\�~B�>�p�)�lF��6E�O�;~8��:�h�DI*����8�P�BH"дԣ�?]ki*+�E��1��s�`�t�*'�>�?.K�-]ąް7>��J �^��>D_	��*98�	���~��\j�L߾��݄���8-�0_�J������NF����yB
����处�%/GY�����q���F~}wf�Xg1��º{���W���aT�������"Ҁ2���Mt�{V�C�j$Y�~9u��q�/�IS���4WYoq�~nt��#��@��F�������
n�bF��\Un��B��HZ3X1�}�6�Q�1W���픃t�#�W�_�̵��
$m470��ID��%(p$3�����[���g�%�3u������m2lW�QV?l�ï�d�6(A��\c5:�=���u�`��xao�|plJ�yL�#�ެ|V�n��>�J��9�"�]f�n��l��㇟Ͻr�������
�Lfѣ0P;0��O,��Dt'�!=)C��F�H�b�,L�c�s6�6�~-�t�R�)}���q�A)�׏h��5������mx���������g��	�ܒ�Q���آWz�cGE#�>����?�!>���&���\�J���|T��ͩ��ׅ\��Ts��D4hw���ܘx_�~y[w��!nVy~�!k��5Q9��4��D���qb�4&0����7��ݽ�B�}?�А�7�a��h��v��8�+�5���lA�~*D{��^�x��gt@�R�$�\��#�3�W9�����@�5W�hx���Yapu�@u�H�m��8�E }���V=R1��C�L�f���3uoJ�~�K�qrŨ`�I#e�L�k�0Σ	[j��{0�KK����<���<)�����2O�r�Z+Qsֻ������Sm[�V�p��vg�'^&@n{M`���/�ء�<q��,���%���1�n/���R������+/IuT����s�j�(kRƑ���&:���Hqp5���P]p��{��[��pM�h,�s1{�8�EqD��=5�S�בKF�3B+���YvQ�B8^���2VUP� ��4�E�A:��6+A9�0�
�%�P*W�7L'B�&ǈ&_bL���S� l���ư�la��7�Ya~��pkB�I (�4�$����Ţ�!48rt���Y\���o�}/cBj-���r)�u��m���o���#�d��1��&.�oK���i��3zO�9�7m�o	�c�2m۫'��x8�iv�ԷM���G�?�#�r��f����s��Ǵ�B��Yh"w�<?f�y�v~8�o�����ʡX����r��G#,�>�%e|�&L�����ޅ7��SP�Rٷ�?I�2�s�Y�AL�N+���?k_�y�$�j�T�
T�kT��O�<Z
�ҏś�q�N��|�h�~As��U݂qn�uj��* ��Ewr����q���Gt(�_�KV���=���Q�K�L���J'���w�e�3!g�	n���<���8���,�a�S�s]�� ��臈x�Dfbn��N�؊L:�~�x�<��*��>����������o�L*�f���K^�Z/j$��-0�9@��"=��vc^�[I~R�w)ZMaR������r�J���t����	��r�9����TĮ�ȓ�x��z!wK�\��Ao���T��Yz�O#�l���L�E̠�<��bs�3�ے��Ȣ�~�J��{�M�H���w���D�i��̕��<��Jlʃ �Z���3f]p�J~�*Ԗ�Ԕ{ȳW��i̲.��f�t�KO���K�ﭢ�Hwd �O�a�4���˦���fCWD��;�����Sb�CBrf�_Ku���5��`���eh�f�g�����_�����X�'H�9߹o�����x�+�Զ��z��.pnu�-3������k�m�^)֯m�4uxک��5�a�'e?�S��Ģir���� lo�-O��0+<(ɮ�ĭ��t����=/���[�9�U�뜰r������g��{����Q��n:/q�u��$mQ�Ť�#D#a�N�����A�`�1�gd��B.)��X�O�Z��Ho���h��f�p�2��bX����u)�!Τ�(G��M*i����(���W�?��}���Ƌ�Յ}�G��mn[�wI[r(HXN��s�f@2�b�D�݉�f*�^�����݋��ʶ(piY�9*�c0k ��?[?���Yk氾�o=�C`�Ti�a�Z`�@�{�o��W�	.8��n�6õ�VVb�xs��۩vh��II]�����\��p��2CH�m�nk�+���� aq2/�o��r�^$��6$c��uѣ^N��Y�q�^�1��u����8�vd�#C�*vb}u��t���8�8�[n�Ikì~�_����T�)��S���4��ͬ���q��%��7A�C�;���vc��>�����X�&�"��	Y\�*��
N}��!�jT�9��T''е��)K-EH37��k��PY���i������N�D�=y������<B��N�0�)���3�ϗ�ɶJ{���)L�s�����B�|B�W���R�u��ʳArFu �-�>�|��O�t��^�O�T������_� ������sZ�uJm��F>dV�4c~mzd��,��:�`##J-T�Z!#���~���ɢD٠dss0�߂zv1���pL
9���#0�)���]�k_�m��s�p���tWH���e�p���F�I����i^X�L_$�F���-V�f�cd�X�]���&��5��7`!��玱3���k�������F�|�ttM焥oJ�s%B=F|?�M��:r�T��u�'3��?�%r�>���hT_;�c[�7�s��F5ҳK>#.齵�_��_�R'G��0�θT��2��ET
��l����o�j�ʼߺ��M����YOԑ4e�]+z\(*���N�=��� @�%}z�:��2�XJ&Zlb8���-�(TZ��ؤ�cw�%I9��| P� q�$�� �P��,���ޡ�ȶR�V��o*n,�z
�����:�b���r�H�Έ��%��HW9��p[xyX���C�k7-��f�>��^Dyîb�d�*��J�N���+�UQ�����c�-��ϩ#` D����]_�]s�fo�Hjqin
?��~!zt* ���C�-�o�V}�6%/���~W��B��^$N�r���20��9]+��˭W�(;)���d0C^�����	8��<!��X�wX�7K��9�= ��	�;����>0��+b�4ǟ���(���Ѝ:.C�|�v�z�� (�s�Y����6�F��aFO�S���b�Z-f�0#�
����9�|6���CTuZ�.G�a����H&��js
<�6�z��p6�_����X�ؚ,$-����Sa�ii5i��)��Wvb=x\�u��Zh��4���.�g(O��*��r���w����O��Qp��Tv���9��i�7�
ʝ����+5���C�Q&)hs���C��/�	�$D�we+s�R����i��	~ö �ˠT�S��4����y���<�n4I,��BI�D�@aZ~t�[��5�$cH� _�+���k*m~S�'�b6�hj��$��@�X����1�VL�&�E7IQ���KE�6�h^�^4gyB�+���@�=�w���I�^Ŭ�F��Q��O��А��W��*o�R��p��j��v��d~��B�.�fr!ji���$�,�.�l�����4�k#����e��g8���m�rƗ�D��Q3yW�YO��W�Y�@���54�=��R����+�uY�j�
�r
=�6 F�����eL=N��0��U�\�R/�hHc��s�d����p�$��D��[����e��f�����w`��z�ǥ���i��������|6�)���ephS��Yb;����/�\e!�wC�I����������+�{��p��:��lF�3�s�:8�|$��G�r��1;v�~�� �n<;�Vy���!S�iߥ"��a��=@��Հѳ6E�P��AoY��Ԯp��x�7�~)��
�},�S��T����Ӱ��~�"#�W����K�����=������V�a����<��
ȁ�suů3����д]���擿���c�.у��l۲�h��E���/=!�<���Qq�ߍѱ=���=����8��D�ã��[o�'�3�mF�����2��۹��C�� �[�tMy���4@"E(�E*qKU����r������])�T�a�CI�Jo���jk��\֗��3G��|����n�8)G��LC�
����s�yC�⁛��g�տ�y�{bǑhT�Ph٧���`\��ٲ�:��Q�!�j�uJ���{/��[��]k��2�[� q,V����X�[Z��;�����|���'`�,<���zXvn��~au���CDEY�Db� Dnq9�Ȼ�f�\Zx��*�G8q�����$�=�pWF  LT��M�WȜ{U��C� 0���0����5��1'b�sz>�lK�C�E�
(5���	��s�W�!�Z�3fIh6������<����W!$��`�a��",ffP#���f������͍l3A�$�(
$f���(>Vr A���,��s��Ԕ�b��E�Ѕ�����k��}�w_����I��9WlR��
��A-;�^%�����H�܈�m�.���YJ�6��1Z�ܺ�u#]Q�r%����C��g3ڼ�H���Ã�8=6�-��ݶ|m)vO����d���q�)O��7��W��b�d�+N[z&��;�h��QNįyi�7~HV0夢�ଯu��H$цS�w�p��0M�g��s�<vt�W�Ȩ���/�J����Ɓ2�^Ӑ>vu.�5y�_p��vX#��N�?��eN��t �3���a�{茊�f�F-!N@f��M�	r�-��3s�M泂2�j��w�Ҥ����6p��g8���=�C�C������Z����X�?꠲�����5�-@�N'�W�&��ą��FKn*y���^:� �dO�zr��)>l^[G�#e$���D�߳	���KP0f��O?���ߙs�<�y�Еby�h[7������.,��l^΁Y@�/��u��
y�)�9���B�6Gèp���K=Ra�E�ph�nn����}�P����P����"AE��J�a8O��y��a�~ᚼ7��0q������Kx�H�$�]��{ۭȼ������UV�Nц@�p�Z����aS&�2f��2�݇�+h
)#�z�'�Q2�F����8����X,?��;n?Mk���j̃{T��o�P��ez��t��yȓ֝"s!8-��6����;|���Ő�N�*T���&M��AG�~N��L썜�y��Rr�+2��¦E��͚�V�:w����y�}O���h�ET�e�r�l�<�$�h�I}�޸��3��d6��T��в�7���YnsN]���u$3�����+9���꺨g��=�ZH�g-��hDm���ډ��jI����4�c��uo�P��J�'�kwm4}pd��̦��-�	���@繨��yƣ�n��nGNN��`�T�9�3���ֺ�xF$�^��3d�&�)i.��t|>!y��F6$��a���]D�|�J���s�W����q��L�ʹ�7q�4��~���Q11J�Q���w)z����&������V�� O֑�L�i�C=�z�1t���/K�Ů�~tizyW���^$��?���M�?��g|@��e���z6����Z�ox�D�eᤅ�9�qa�����`il�с�{�*`���S���B��a̐fb�V�e�[
N���th{��H)��ҷL��<ݔ�v�m� �P�s{`q��/�o���<������-�S�P���̰d��ʡp)F�N�5�L@U�A2d?]Ǵ�^'���3��}��Uy�sT@g�>	Ent�;��S�k�8�|n�펝��}�2� ��9G��dU�|��l2�:c��{��Nv�r2~a�s\���KCY�r�g���e0yz[$��&(��h=BH�����_�_�<7̾�w�N/��t�gc�� �R-��i���:���������=�ol��h���w�ّ���O!�����~�����&��$��2>�<#������9Ἧ�� �5��(&�����8�Za�Dm��;��V�PᯖV���cWP�`~������wc�]�^�:$�[���B��h�}U�q���N��gZ7Lٔ:r�2�4��Nwt�'�9P�*gK�(�AK�-�)�Ƥ�HF~p'�ps������L�u'-���}��-xƣ��ѥnM/	7�
����>@�3����&�}[R��T���ϚG�9�@W�7����c�\�#�6�:�'����|��A�������m�u?�X[y�'�GT"���;&
��`|�J�v	#y���J&�ݩ�J��Q�v9�~oq��*���HY?�-�dwl^�?Ӊ���W5���S�b�j�:��*#���a[�4���a�.�~�*�2�ެ�c}W�㢵r����"gh�0�1"´��t��t���M��<�m�,"̂�5�@%`h�>f/d��as��1E{�~���e����Q"�U�����!k!C �iP1�m�x�t%����q�J���N��+�x�ﮱ�;�����zafX��S��e�5��7<�!����%U��虫����RTq��e_�YЙ>'%;��{�/����i�jK15�{���ľ� ]��������-A���^R�~����v�Y�����pt���m���ש���!�(D�lpg�C��(�f�-�v'5*f�)�y�~��y���I�E��I�ʰ|���5�`��o�G�t��!%
" �׎���eA�{x%C�����gGZ�;hpv�䎩l�� 66O	K�4����5��Z?��;,�����n=�����t��C
kD�֗�P��=�%���L#�/�g.���)�;�x�ق)�U0'q
����zG�[~J�ne�J�9	&���s���7�wip���/M�v��Q�wn3���P���XK�X���XN��
���o=S��Sc�㿜xr��܏��*M���9$�^�5�)�4}<�_��R��� �mD�ͨg�H��\�@ێ:B5?���a�q��[��kr�{"�ۅΜQa��3���3â���x!A���9]����p^2��lҳ[Cm�H+�tV���ߋи-~l�x6t 1-����	�y/�e��#��L�/ȼ^��ʞ;�8��.$fb�$��wΖu6E3p9�2:���[��}�`p�Oun��k��^|��ۥ�h�� ������'v��5�I�+�y�]:��8�[��U�0��RC%ҙ�H>�x���/Ҝe��� wh���i6�;*	���:����{�I-�P�'���I��T��yV)����T:������IO�Ar�}o8�T�1L��*�,}�E�������Dj]�_Z�����G;H+.���h�}�~��^$�����Cp��Aϳ��*�y��e��7�X��u%���۾A`!~��C��By��n�_�CAn/�����J��W�����N8��s)�2�6Ƈ��na^]Y�Ē��J�쌿��S8)k�I=r��σ2�.+Z��BMpi�@�:�w�RH�Y�BD����O��~�W�l�z�WS��DAM���Ok���͉J!��~�κ��B�W����jm��7a)g���DT�Ŷ/�k�@�m3�OD���1ߊ1p=�0�Ρ�x�+^��n^A5�(S�4�$8e��od3��c�D]zi�n���<�t#�9�陕�Ew�L�7���}jq<KN'�Yy�ӯ���	GvkE4�2� ����<f_
�[��x���$�w�2w�#U�+�3E���K� �d�D�v���Y��c�͈�7E��<�>ci}�[v�N���,A~iS��dt��M��a�������T���1��]�i/�je�*�x�. XO����/!����QI��L�)S>�粞+,�[���f6X z��Ղ���K>g.���=����E(����cbPŇfh@,ݝ����h�B/��������y���h�K�D���h!��gJ���)���F�,�\�KD��j*���yZ�.j�������nt��An��ԧ�n>ȾKUօ�*e�6���
�Zwܣ(p����N�6���M��寀�*�T�F&���%nƲgCԸ���H��$�}����il�2�$?��d-m�MC/�������П�LR�d	E���~�n#]3��G�Dy`L��?�)ߏ�0��5.��7f���%}Sq5�*�n_�����Mwī~}z�3�� n�l���a�J�yspS,Ꜣ�-b�H$-��7��#Ym������)3�~�[/l9vHW�\���F�V
3�a&��1��m�Ʃ�xauh"a��}���[#����'��K�kA�ڐ���o�,=]�����rQe��#��Z�ω|г�2)�@�{�i�8���i�0A�s�G�:Lz-j�Y'��%I���G�\�)V*>�pL�^gے�A@%��2Ů�UԷM>n��mƋ��l|ac>�N�n�~ڞ�����З![����GK;�
���Z�S��_�>U���8${�w���J=��ݼ���c�t�p���W��'K�0�vv�/��M���� $�U��#3E�MfO�,]i)	�
�X:61��v���Y���b�]�|ͨ?X���gzq�<�h�س�NST�ԣ���9�師�?f!�%��8��x�^�G��ƅv����ߔ
!���*��d�4d�|<ڐ���F(	�c<�o�G�)Nx�Nȣ5�`?�FSCլb�*���R ���?�Jã�LV+��'���ק�ǖ�k�r`D����h&���2"��&��3��E��6�g�ګ��o�)@��(_k\����2�6ˊ�H��8F������j�P|�#��������C��Mg즆w�������Ԓ��J�E�D�neXz���	hE/��cG{�~H�m��"U�t[�꾞�S�!
��V��{H�l�]<�>>��ϔ�T0�� ^��[P�"�;*^.����O:�	�_�ʴ�eϑ�` iB
�5�7�����?���e��L�,6RxVU�%���ތ}u}l����Q���F�9˺��7�u�"�g3e�ҿ��68����y�۟kʂS)�:�{xj{�C�jux��)�͈s��^'�D1h�f	�
%�a��EXsEm=ʟ�
^W�%�O�m�&�V�"N>(���EK70�v�+�@S�|^IH�1�\�Pp��T���̍@����@�`s�O�CMq$�9�`ҪM"ءl��g�Ƶ1a��u�_j�5�r	��fɇ��묹<l�P��'[��5(���Ԡ��=�y|?p/kCF�Z�MX��0�<R�w���G�"��;�m�Wɯ
q"�&&��Kw9�DI�,ƶ��X�<��K�P�ŗ�Q�%��>��@�������+�@nɟ�y����Fq#���_�M?L���%�@9Wi��K'w�)Xs����p_��Ez�iV2V!!�����v�Ӫi�� 9��C7�mҤM׋�5�4�s�2��c�P�9�F�9�Rri$�#��g�e�z���Z�*��PV
��ƚ�ո�u���'��Op0��!��)�Mq+�9��/��$i�cڇ1� �7U�%LĢT �>���݀��$e�K.8l�=�aI�"CC�P�\���ujx�4��8Ǵ}{�~��;S����+fAݕ���h6��Ϩ����-�%��U)��
VaX���̳�4 ,�Oh�<����Ս��YW�B���-rO�|��A�']�S�Hmm�\���vD��j��H5�+��JQ&�|�";��lQ[úE�?�i�ƎV����uc����6�s��	Ȑf_w�"rA����ؗ��#��r�Z��vp+9��i����I(.:�
GC�w����_d~������#�#fa�.���Wqz���C�X�M0�i9[��I��o2Ǆ,�Q��6#ϯ ͛�K`�MW%���P���v;�{����
2H�r��逌�R`�4 ��c0�]�@�v�hb�)+@��X�K0�rniE=�^&]$��#uv)Ts�8�&��4��c(�N��t9�5��*��9��ǻ�3"Dྲྀ���}w\��],�Fr��9x}�隑ѐ���L�(��� N=�R��$pY�>_�Ÿ�$=��Z�OҾ��i>Zal{ݱ+�^�2�pnD1���̾�EAv�J�}?Ch~��?f����������L_
bQvXA���%������+���P5^�=0C� ��#�2��GXU�oY^��j	�Ur�N�t���ߧ�[ky[0�s�5��`r�h��Zk��Sp$N0�3-w�!4�	�"$A ���(�
ҟGsN��?��#�1�]��B=�f�Ӣw۹��P`6>8�@#��%���N�K���;ɢ%�Gv�)�P4n����i�5�c�P+.��
����a�j����1eL�9�2���0��C'��P4��q�{�ym��b�YyM�(���)A�K��+u�7��Z� ������E���P��2-�2MH�6m]��-P�b]��?�z<,'Vw����&�1���ç�h!�%���)]��ώ�W{�k�	=i	,��˟@�sʓ�~D4�h�4M��QMy<�⢴���79D�΄���� �,um�/�����|����Ya����"h���da�Z �!]l�|���]ԔH��*��fG�	�7;���~r��ST���R�w�٥�Q�n��b�d���X r(�j~+����� g'�"jW���d�qr�	[9!���3E�R��]�g�?0���q���U�(� ����5���-���L%��Ѹkt�:�4~3��}��hl������Q���ї�u	�P��hB#"�c=�<'F��_"l���^����Џ<��G�A�U(��]��S��VF�Z9�n�Q�q�{�����t�D����s�I�?4��$���t�$�{�'R��d��je�]�3@�������"BP��	2�9-�,���z�� x�,�RhX)*DZ7���`�;��|�_p��8+����9�,me�R�a��z|���W(U��>���~=�͞�EPk�Sb�J��^���6�V���mB�|�ͯ�) ��|�W�'��j���,d1ڣ�B@:΍���N���,F̼�K۠#@ b~�ػ�+O��t�{�o+�8\7���^���Q�.S[4"�>M���3W�T_��
�>CL�iO��,�y�*��=y���vFsO6�EG-I�,@F_�w�u�rҬ>�%�w�������Ź��|Q�YM�y��n/�iAϣ��HȒ��5uY-seD����)jP���.���8�`��]��K+}-_�9x��v4B��Փ�n���9=�ȡ�Qmˍ�B���)��n��������Wr��b�&���rE�g-�|���0�r$�PH�~Z&���-Ź�f�.Q�b����3�N�u�V�b��ϟyE�r:�`�M�Y�s&��*�6��9i^Cm���AVB~�t-�Y��OړL�稓�XZr|���Q�|y
̀����)�����>V�yo��܌'�.����!�1ʍ����os�)��3=��=jJ�{�ұ�aK�G*6-f�X���j=�u�Qhm0� j���n��)D�.�u- a�֮�k����Q�b��2���cd�?ɻU�����ß��tE�4�%���1ؒrMF̟��;��c�	���2V�u�a�h���>M�c�L4m�;���V�죩���w�!$��p*��7_�Va#��K>a�(�����z��Fͺq�F�A8j����\Rh�mx��V`I���G5�:����z�-��2;�$b��a+���-��Hh�dҐ6U�Z�ۅ�8�!07���7�r���$m��%�����2�|�Y��Sfz
ٹ��b�2;�5v9�NBx�66�ݧ�E ��_oZ�P��(�kF	ۘ�݉����k�6�"��Gs�Y]Y�hK��^��o}�:�/�`�>���/lWB����n�P$��B�g�q�
��|/�9`����F�^K�p���M���k��83m��1��#�^��2�b�rHF�>0�	��{����X�������\�h�up��<C�^���Y�RC���պ��1���X��G�����g��[���F�J,u$2|����������$��\�]�*�=�*VX�5��ch[~?������p�!}�)5W8�*���t�� �Jf�%&<Х�RRs(:��ۛ&\��Ī�.k!�{�%��q��e,�0��A3�tu���"`��
Qr�!擄{�ϘW����:\�U�\��%�]��[P&̇�q�}���j�r\� ��đwA�\�����-�)L��Gn_b;&!I���h�P��aK���w���݈�`����u�Nٱ�Ѝ���#l���h�	����8�]��at@�<��r4�%����/��is�s]S�*�96���Y���-�5����1,��l^�z�����Ѝ�.�"�v*5��вnlO�&ej����8sT\狠��v���w��+�7��9* ����$�\���̐})A�*d�a��6x�B����}v����fl�'���/^3�l��u{�0C�2�SK�� 0�#�04����ޫ��~�i3Rr#�
'~?
Vf�d6�9�F5V��]D�1���U���
��*�o�"���ǎ?��Rܕg^����]�qa�'$iE]p�8��H ���u� h/.4�eE6L+����0*:��������y��A��vzyZLz�c��4\�OjC�v(��a-w��	��yh�in���T�*i�  8S<�	 $~R��J�s7�v���ԟ�8�,ج��D�����u��D���/:�y���NH��!tAe�_T�G�ܵZ�.�W?mHH��>{m�D�v���Kab�FV+�ev��ᖲ��C���<�
Ks��n��R5#�EԞQ7Hۤ���od���fOz`�<)wO*Ò�d�"L���Ih5�#�f�iH� �̈́QS�����,��+��f�9���CO�q`��CM�d����"�_ݹ��bZ���'�f�v��[�v�V�R;��.��s�eE��R�E	�����G����=@�����x��j��Y�I�Z�N��S��w-yZLt�ȥ�*d�G�~&���2��
c�G��^/�S��<�eŞ�rI�T��Z���e���f\�%�W�#�cN\hS�,ޞ�/{}��ƛ���ס*��I���&�!i��E�j�!�H�}�2�q*�(h�DT���\ހ�^l&BA(=��a*(�]�?P�%�m!���O�=�F%��d���R�GbV!�Cz(��=��}��.��S�����X;4�t4 m�Od��Q�}��Q�F��X����}���"��/�'����4�������EPo��UK���۷%d��4 R��(s��W�ys/��x#��Е�Ȟi�ADW������>ŒY���҅U�������	:QcX� d����l+�ǁ(ph���(Z�`�`���sG��	��J�
����r��h�k���Ӆ/�C	�Lr�ժ�э��N��H�h-	ayW[f�㪀D`�o!�� �xu�T?��a��@�{?ZV,���*� �!�l�`\��),����qͿY"��#d����.sjaz��<�7�|�0�Agv
�l2o��Ũ�E��B':�,zLpn�YW��*�*�
Ϸz;@�Ɣ�`�0����Z��������r��lj45�<�0�=�)�1��m�ET�Y���5"m{���l���Q�%��+�� �Q�7u���J����g�K4�h.���~�	�%%����pګ���P)H� Y�%�b�����aW��"<-��/9�Т���{nr����  |�� �Ɏ)�?K
�o�^M���(b��!�13q��5��I}־س�`C���ֻ�~E{,���9C)C�J�kM9����+�g��kKs-9|¿L�������a� �T�+�%	�LjK<�Y� �����6[��΅�
��*beo��.�OQ�����H)�n�d�aJq�������i� ����zqu�������7��k�p<��~����NيJe����ld������W���1�L0@�M��!� �d.`=KZCڷ��J8�*�3�"0�����e�c�b��3Ѐ��P���a�=����'�xm��uU�8����6n�g���+�Nk����1(�ۻ�
gD?}p~�(GX�Abw���Fm�E%�?��"��TJw����i%�	g���H�t����/G���.�����r���Zv,����R2B0��ֹ����_� ����X�g丒;e�\O�[�`�ݡJA���r��4;ha�<����o2�;�{�?�V1F��jE��Y�Ѳ�3�0���Q���V�q�W����a����s���;�E��uŘyGf��M�O��N�[DG�í��� �S5���o�fֈ�0�i.�:ɽ@;Q��ךh&<�KmKQ�}��M�9�[��Y0��I�*'�Ӹ2*��:�z3��~��Q���`eU*eC�c��x7�:�����:�B�����j?d�
�0c�(���Z��7�y��M�"�"q\{S*��X��t,�+Pk^�J�F�.<��I~��6�v�w����d�����}��l刁�-	��jH���
S��E����~6��h{�Y��q���w=��,�Ks	Y��v�.?��0�-$��uI�H��=��L�j����T�#}��O7�撢M���Af>���.Oa;��FAp}K�V~���\B�o�������c���<�r��WE��2��|�o|��X��+�v��mk,�GձSe��h)�2��5�Q���T���(\�R��>vB�����y���J����xq�j�E�%ȓ4��;�!W>��������'�?c��l�U,�}���qckH���(U��'0;i?��Q�����oe��f&9E��y�^X�0I* �)�+"� #���D=C����%�\'�ź�(����X�GS�˾%LJt�W�U��^�g�������/�F[�gx�꽥S� ����N�Q��)��(*^[C}��R�{���ϴd��bۥC/i����n�I)\||��ǽn�x���b/�&�.��0��e����~2�yi W���E�����������&a�\�蠌W�O��"}�`�����!K������������ �W�[V��o�E�m��1��,���r��M�}���c�(�\����a��R��zYOR�b���
�5�8���c? �u��r~,���7dS+�ׯ�za�C�q�\lH����.������d�����Ҙ��&�dgp�2�7�IZ'�qJ��Be?�"�� i��&�dC��gB1�/$�<�i@z`�c$���G�<�ɫ�-��ɕ�܉��a���H�\@[ϼ� a���o�Vr��f���<ݥ5#���:WC2C�\b)d��G'C����|H�̛ R��l͟����6D*I����&���I0F����	D��'�2#�X�(�f!����åAh��Lf�{Q�l,��Gp��d���E����4##��򇧚w��Y������(�m։��J>��kY�_t��r�H�)�+�4�~~Y�������C:��2>�x��	��,��ۙ��Z��ؚl�����pOv�0�IeG���A������(�6����@'�J�0�Z]�̃yb���\�d�j���?���c�����蚅�ɥ.hC/�#8����Ԓ���7�gQ�:�kg���pNO2)�S�wbF�w��Y�5���|�;^��^����ΝL�=c�7Kώ�@:G�=�AOC%��a�1H	"�~��lF'F���g��������������a�y��:4S�����D�H�]�w��%nHF�Ҽ��8���*
��e�a���(�;&�"@���[v�;�-u�oib_|S�>V�vD�a�fE���Q2}�C\���IFa3������?>C�O�<gE���{��l����r&#�O�m���ru�nL4B9���))�qZ���u�Z��Z@��a�©]l����Œ%���I%T��ˁrʲ�=u=l6~Ú�1;��lSە�KC3��}�e�W�4 ��"���=.�s��5�~���N*�>��s*]�4G�=s�á~j.�.sQ>��qN�-n��f���~�5����dt$�G �Q�ɐ%��2�}P옪�Q�*[K))�.�����f�+��*��P>�3�Ѷz
�+���_��t��2wܞ:�ܓӽ	�쮌帨OcBG���
�I��`����]a�#ɲ���[E_o�]�m����Q�^g�àJ�g���%X9���i��H�ע��u� �a#�X3DAO�|�g�ٛF���9�}ΉW�hj� %0��wκ+]�i)�k�8W�?HRo��� ��%�ێ3Y����jh�t!�a �{����c}�ݪ	��pr�%�-�N�}�ЍdYZL��ۿ	J�}`j�@f^	�K���:>�=�5wK�]h֧��mt�tRh����͝�����Fh��f�W.�
���p�oˡ 	�-� i2|�`�괞ko��/J��1?z�͓w��ymO���]�PP,6]�BX�ǘ�
@"����W9C9�[Z�W�.Z?_"�0��M�O߹����Ù<f����QB��A��ws��&���5��"�s�	Y�%|�*�k<�z�0���{�p����v����E�˯3U7*������t�e�	�y��n���i"���>�e),�K�S(�;A,C�mAbw#��C7ļX���h��zи��a�6�t�:@�{����L��0�6-v�<� J�'�Pje,�y��|�%����6�+�w97{�o�.9!��-�5�,�O�Wr z'�;��9Wy���v�q�j�������63�T� ���&�cp��1�5���F(4�JW+��U�o<��l�
w8?��_�n5V����
Aګ͉�w�*�������Y��C.*��$�q�&�J�^1"�U'�W1{�s�`��ib�O'�S�+�q�`v:\����s�C��DVo>x~B������x��}���g�qP���I´aXd�۸Ѣ���װ��=Ҫ���̱��!3���ݳ]�N�ɕ�8��L�s)ˉ��o!��<���ж�)�To!�߶y�|���|��E42�	���%���~�(Q��/�br��2���$�Ѣ� ��zx��k����X��+Ť�:���痃����7�cY�J���LB��k���˕2�ҟQΉ�erH�i@�8w� j21�\)�Vfl���4�v�7ۇ4�G���{WV�ᬨ���v�ŏ���eG�u Q������;�CGN�� ��.��5�|�o)0�c�!hvM�j��v���].�k���y7�}��?�w6�_�lY�|y`� ��b��?,�O ��1�*�w"7�;!z<���l�Ң�o���T�M�jD�	(ڢF��sZc��b v�@���K;˵ �+ɔ�-Ue� ���pz�~ˊ�m'#HH0_�Pc��W��S�ʁkE�G��/ý��D� f=p��<����RT ��o@�Lr0�*ݘł���
�$o�N7���y��v�,�PL^�n-Dou ՗��AG�O��M��'f�е[Q���0Ǡ4��+�EQ�O�%�\� 6��\�Д;H�K��#K+���`�&3!	�Gž�#7L�p����^\b�İu���\�<H����zؒɴ
VE�ϰ�C�9�2���d�YP�XX�!oW��J��m9�p-��d�}$���f���5_Ty�A����~� ס�&�»#�#�3gc���ҕ����t�~g�'8�
��|���D�t��|wLYzuT�NW���O���E�3E(Tp�Mzш��P�Cܲ��(d��|(��	5�͸�:���o��h�8���-�yE�t�c�eO���Y:ջ�+�^�����W\�+F� L���U��N7�n�B��?�����Y�W��:j�Q��9m���dVu��*�ݿL+��%��q26��~sL��I*��w(�{;�������v���Y��(�-(���b)�޵\�y󥟥�"qԬ5���b�8�����$$�i���ep�Q�ON9:�6�g���Qggv^�`Q�v@v��lڦfC�Nay��SG���K��p�$���ǩt�[��.;����3��[�H ON��#�2eu��u�mt�8�!9ʒ'>@����_x�o�q��"[�{9)f8,���u33ɗ^������l>��ӻTHi��sca�-�����ӷ���nġ1J��>����>�n4��c��@Q�خ>dW�?����"�w��S�/�4$X/s҅v ���1����uv��2J�oN�5��P���;���O#~OŇS��w�O�X����J�LɈ��^y��#ˡ����^�4 [A�!,���؜T8v�㚶v��U��L:��� ��Э�ɷF4V7����ƴp�jF�|��-�9�<�&�\}�ø�?�CS�wJ:ε�c��gV,x�p}p������oIM��7�5f�j�=�ـG���?O�/���+�:Tn�-�Y0Zx������|"C���h�Y�.���ni�6%|6�r�K��зxR�4����]��2���z�D_�ې���1���<B��~�d�1��ߞ�7&s!E�����q/��<��u������JV�!���#z-��90�7K����+��9����vATt���Z��� <�#��,�O�K�̛?�B+/W2'f��真�X�_-�M��O�zHL�7��n��g`�8��3F�ߛ
x���1OZCd!g�5�8%��;�~��?��$��t�[W��į��������V!&��x{�Y�8��ڛM'a��3Dy@�]WU�A�V�#��w�B����kM+�6���S��N�M9����N�(#&�3\�ؐ^7a����� Q������S�&Ӂ-Mn��� O�9��B@������pf?C~�@K�qY���:��D ��1)6Qn���bc��g�����	��N�����Pmy)��×y(sf���?z�\=g\��>�N�����:�������������F�.��7���T���(���C���`�wUx�%Y����N,2��!8/��A�N�~���?�*��4|Wm�vw��mN��c��FF�?.?�F���p��"I�1��ݎ[Pm���W�u��*����ک��5$&�0�r ���Z�nJ���:�. w-/�|uͦc	��|\���׬��dPn����������-��G5���oT�����F��М,XW*��wHH`'�@�vI/r�L<ǒ 3E���
o��F#\�i��%�^�I�Ka�w]�0J�S��\NDk�Ψr�8���
��������fG��������:z�Q���,�F��1�f�_"�$rS[�.�h�f2��Yy�ʽ���QiZ�0�n���	�(��,̧�v�sf��m�����Cw���&�8a�WX�O;*Iwb�S��Z11P	��JR��*&8���v��E�F5�/�5��.�y)K���8m��>��R��nL�. �Z���
1��螂O$~�m	��x�Yg��������{�1u}�5A��(n�j�ox�ك�O�t�Т|�-j-R�/N	�X{��X�,���r�����6Y�Au3��p�! �DP7�-�&4����/�����j��x|�J��l���vGkw��k�xZ݈�y�oe��� ��glx
29����l9R�g����{��ەqN��R���ip�b�@��z�V�ε�I8��M�i�.�C~P�^���
g@O] ����d�ݑ;��ZL�y���v)�C};ս��2(�ҫ�]&���U�\��/���������1��ԌZ_Л�s*����*���I���2A�����\�r0o�j���kF��$"\��}>č�˜�*r��uǜ�����SZ�VB�+:��^���3����:[@oJ&4�O#�8����-)yQ0��2�z�:3��$��/��qo,�FD������̗v�ÜWM�&3��ҏI�n]��n^q̪���pu��?	��I�"��;�fe��ܠ����C��)��g�6���=�����&�����O�����)g+� �q���l8�[�%;Q����0�:M�e�Gi�1S��(����=˽\D��@��y���Z�o8������1A��O2����p"�@�gf�Lw��/�~���~vH
ƿ�@�f�eɺ���t4���v@���Z��7�u~�����RM�L�����q�8����L�9��k>h:�F�ۓ9�9"JS��|m�)����h��m��f��Ǭ"�����˰���� OF>鿈).�����y�Jv>)ᧁG��z���+����q�]���u ns`A�gCX,K}΃QF
�@�Ϭ�̻-o��V���!�j<�� ���i&�¿�r�[M��pJ���/&
x�ٔ,��1V}�����ufҤ�b�Y�@���}m��:;c���ͪbqh@���DͭP�-��� ���2�H�)�����+�|�>��gG�~YŇ�QIuN�H;����JW$O+sY�<�E�@�}�a�?c��j~����jDl��4�Ս}
����� �)�ʬo�G��u F$�\^ri_�~\$q�i�?�OTqP����+��+��@"G���Iy�(�#u��~��$�5Vb^�~��%������ǭp0<�ʫ!;7}CJ��w[���y���XN0��M���76��c^l�e��y��f�J-�"�=�09l.��7(�����	͡\)��
|�M����]L}�/���"z@\��� �T{l�~6LG�,�(��);�>��dTe7��$|X){u�<����i��;�\���Ὼ��ZM�1[�����|�9`Y��z������%<��2�Ճ_C, w�) ��|O(�e��>րΗg�"� �#�!=k�B��>"c�~�!�v�`�c�v e�,���H(���3����M���q˨�4�;�R�&~auQn�a��aOTq�0M�9���̆0 ��Z���13ӥnT�y�Y�Uʆ꭮���/��sK�_��Y�������bWdG��L��K}��R!�L�
m֋�-��~y�_r[���ؖ��>�и=�v��aE{WM,������)����!yPa&6�rӮ�q:!ݭ���|��@2��p(��8|#:�z��s�*���dQ۫DN+ƴ�Pzk��۠`����cd�Z�J�vfp��(�������O��+�M0g��,j��\ǟ��K�.,��6����;w��-�f���)���]��^�9!|��M�`��Ǫ���;'i����e�������`��n�"�2�
������c�-F
��Ҷ����l���"��:eX�K햊��,��,陙�4�k�	�9)i�d4̈�I�lv��3pk�C����~�ۑ#բ�(�Z���}<*ɹ&�Vs8h�?[��`�Cg!���j��ʃ묄���J]%�O�"�~@qȚ�I3���.�]��K��.0n�
MH�� Vb _�+�7���,1 �6"���f�2��7q��W�_h'��;T�]���K�ce�=��kc�kߡ�NA�BP��)e#�&�>���w�uHL�x�W�鬬V�^�L 'y���d=��8ΗsLm��[de����m��ӷpd�������Ӥ�T�H��[��W�+:�8��%L��Ty�N��;� ����
�އ�uދ뿩2�0�&���a<����׹5:�+b���N�]��_�QO�ھC3�W[N[�Fa��<�]{�V����>`����;���
�4�`��3ԕ��� �=f[y��e�'�@�zh����1��x��G��^�xd�9�H-@)�����������O�A��L���,�j�2����4}|���?�'CFo�ܥOk�n�:�N�Z��x^�G̸D%ɘ"0�d�i�8Ĵ���fpPm���>�%&�u`p{��l
�2w��[S�/���|i׷��X��fM�������G�+w��y��7��4G5�I&�kcS��$Sk������v�_t��|}�rq���O��^N�]z���}�!�Q���u���?�k��/Ou}�"R|�c2��z���y��U�,�4`Y����g�d�+�<�~V����8�ֹvAx!N��v���;�;��h����b+�o��8+�z`{!,�ˮgg�� 65��"�Pj��J=x�e��׽�n�$Z1�A
3��i4^��%^A$�Z'}�^oi��m��}o��(\9>���1a�'ZO0π:FTƇix�\my4��^���81	�Er[8F ��������x"�ˎ�k7ƥx,�������tS��WGj �׵H�M�@�>#�ю=��@�f����Sk�*d�0�4�?���6��5X[A��܄��x�M��gR��
����ͽލ�6�!�2J�d�n����ՋA���{\�q=�����*�҃׳�.��2|���M2�Eó�_n�?-\!�1�3|���!Zt-E�v)f:ń#��M	d�<.�+]�pZgad�7�R�⌿�a��~��mQ_v�#���ϊ���Pq�<�l?�~A�߭:����,}��!("j�7�J���N��͌?�[�J��Q4#�u�܆����H]R�q676^~ ��I"J</3jahQ��s�[�R6�?s].U�8�
 ���C��j�����e���h=Rv�#�=�����U���!�� 6�B��+�-��Q�Hq��	��z��/�7$��[Nf���������s�} �J5�[bl�\`zo��tV+�<W�Qҟ�3/��_4,�ǳV������ J���G�,qU�qt5����[TW=�e����f�6!x��1,���J�v�¯>�5s�	��pe� ���z�����0�8"#�<��W1�1�Q�^b>�w��m����K���4v32�16�?fUu��V�uN��=jl}Ho�)e/�o�#m�!m�Ac0� ]�~���"�gX����_*�����6��f6��Zϴ�B�j͇O@�B�
�l�WLz�0������po���(hG}�~5�m�U%����;�ښ�TI)�Ȏ�Z���xgŶ���Ҝ��g;��2Nf���I������X�u�'{���c�!R�@��*y��
X52I�j��8��P¤�+BP5�6���L�K8�kXV����5tD���Iql<����*�ұ�)H0�:*t	Z�Nf_�{��u?L�����1�ł?.S�\i��-��{��i)�Gjx>.�����@����=����o�.R������֛dQ�I7�����?��ʭ�ʯiJBB̸8dY�}ǥՙ��(��'����84qa�-�����[	���?�?w���w�.�w���R]�)C��
GK�� �a�E�:��]:����U�b��:��V�-������;����3�(��0�����:���E�؛"���h�N	���ʯͺgr%���L�>�����E��[�#yW��:����X@U0���'���AHx�
A�O���F��/#��}X34�� �YD��!3'�%R��'���"�Ѧ��Qʰ�5F>w�yۤ{�+Ih��L�sk&w�6i�i�y�}�ƢR��P���r��ɰ A��z�́�zB��ѿ�
�j�:�4�Շ���\`5'�^��w5'�|�㫇�Bf�
�+�B�r�0����D8��h�ߧ������Hc��QL��\�1��c� ���0TΏ��b�\1
s��:ߐ�= �/��@���z��� G����N�r�$�z�qƀ�:J���_�1���ʛS9' sd�n�+������l1Eղ���d~�����	�G�]��#gx0y�e���zz]��
_�!}(#�"Aϕ�1����Ѿ���X����6z����]^>��M��\����Nhw!)_�K�DN��erzfv��}���DkIя	�w��Tc`���-Z^+����31#+��6�B2�<��N�W�y���[�;	_#P(ou7-,��� �m��h7�H�Va�x	�Xi/c%��l��LA�
�I=:y�g3A�g1�4ϡ��v7��񈂄�N�>�p>B���~}��pB2r��wS6�+޴B,�؎U���T$��k����<n=0[T?�Ѳ�����~��+|o�PM.��%Ut���iE�V�aW $JLͪƬ^�_��#�Ĥ�[N�E`2rۼ!��}*�O�*W��_�M<|S��St֝?�!�����[z$���o�>#����B��лҾ�s�)��ǘ�H��
�4���U�0z���)F>a�M�>�́��&H+�2e���n�o�l.>d6l5�������e�n��z�"#R����l"�FerΏS<�<���@cA��AD�x�T�]$O��褸��HZ��]����%����s�e����#R���d����?T������<�q����o��K����CA����(�Z�h���h�]��xοC?�t�c޶B������Y��*?W��u4���#'K�cYg��1��=	�yy��n�I<+��	p�bi�on�h��x��ۍ����~���}����7���_���Ao9�\��::n�Ҷ�0�|/}n<l�e1l$4�a�y�� ��0?P;���/4��z���h�}p�p��|U�86�#��� ˈ�ݡ�O|�:�vbF�1�)lqw��BIjY)G�L�i�� Y���X��Z�"�t�M�>ީ�EcrP����m㚴`��czၧ��N���)��!q�/|lT�j��Nada���,

,@�����(��`g�yMD��5Q;��g�2׉آ} 7J۩0�6ڝ��)�e�*矘1�o��N��&�ˬ)e� �J6��!~�^����y��Y���?]E9�<� {�U ��U[p������p�	�~6�����W](�V)���g\X�`#��E3o\����k�G!���ܖ��;�v?���|A�?��@ �|Nc	?�`3ސs]�tz�]
��p�ԅ�UB����?1��i�Ռ��N�PB��v�󀥤�N���T����;�l�j��нQ�>�f�0�N�Tŝ��a,�%$����C4���k<���o���3�Ϥ�k�vO߾�5�U�GH�$utA�Ui>����'�D����c�����ى��\���+wnn���-i�E'����V8��__�wbbp2��o�	���!y8��y�em�)�۝��5���\�D�
.���!��e,��z�$ɟ}��t}VtT-���N��W����`_>Z
K��5����}�?�z^��s�q��5��!ʱv"fnd����#d�Фx��G9;�S��+,h��n��H9b"���� ���{ˊ�	�a�_@߹c��|e�["'�Di���N5��Φ�e�Ɍ���M���+���N�"�g1cm�y�1E�����'0�]�8&�B,���T��t������@��Ι����!qo�0l9� B�Ƃ�p�5�(]i��)Vz)���<9�zp�I�	�f���F5����+��MPf�1<ߦ)�DO1`�(P�A���>G� _�נ#\���
f���/lܟ���B�Ո�����F�As��IG��+
_�{���KU[�&5�Z�#�)���^X/���z�ֻ3X�{;���� ��U�o�A|�v	�~ƤR����CnD1j��|gT��԰�
��~�rܬ�Y����6�ft����d;W�� ��`��(�I�H����U�K�]�zT�;�\��* 2Ԯ{�{lߊ/+�2J�^,���y<]�9�nG�3W�p^'������ �m.�x�mrk����d��(��Ob�����g��V�z�.�֑65.U�.(p��ȝ�`
�J�K=��|nZ��ް߽�(��G�~wD�:N�$Æ�0Q*�^���Rj|��pw-B�J41�_����I+:��z&48� 0�ڗ�tZ{a��2I��Z����|>�M2�2�p�|�A,AqO�Y��'-�W٨c0^Caϳ�D &�缠�+�8��/  �?*/2.�6�q�g��b�6I�	m�b_{�T�?�>���*b���U,[+{�~_��\h�����c�E��y3�5� z�۴��`�K����;������O��� UA��s#�榏�ϟ��Gύ��4)ς�y�`@?tޣ�PZR��V�����^������&*e��e�K��_�N�X�Ed
Q]r�Kj}�|��\��ȸ������Zs7z�ާB�&X�նD��>র1YS[��*{�bUhnR�hB��h��V8�J^�4{.;�MFjZ8t��:/G�Ƥ�  j�}>��d�C𳁓�z��9�HxDy�g�,�`��Q��b�����L�8�����uI��j٦�"t���"�����9��%ƌq�ثz	�07��W�V&���4�2�	^]�����b>K�2Wk= ��F�f�I�MB�$s�k�ȉ`�q ���G:VU��`��ݦ�g��'r�������Y�af��p�x�i��x�:�Y�ī��TZ�X9��ꦇ����ꌫ	��S$_��3���Op�s����J,4rT��.�PLj���	�,�LhA˯���Ƀ���_^'��M����8���d��6|��ڙv���ʳ���fz��M��)���X�M�~x���ǀ�ܫ�Â��jKul��NG�5.��m+�8ʁ���v������J���}:�߲x�5J�c�����x��WW�CL�{GнClv�T<���Ķx�m���E���Ek��9��1� f����J�Z_�X`�-���Y��E�������/'�@6��]�#)x���O�{y��ns�L�f�z)�a��F	�Bh�$>��;,Wa�2�T��m��_�l`�/��+�&�3�3B�.�
0']V�e������1�� #d����wG�P�Bn����d�wńE��j�����;ڟ��#�:������`�����D�RM�����gd[�h"zQ�{A����AI�i$��-�'�,sd�Y�;z*�탶E��.TW,��e*�W�}��B�����&��i�L���-#?��"�߷�����	;�l�M[|�]ϩ'sKc�z���	=p�MCy���h����z��<�Ou��zL��q���JX��r_����֞v�ۯV�w��̾�e�`�\�F��ڹ���0�o�@�����a�pm� �|�9Q������p�	��YbH��H����'zX�ձ�~4��Qh�y͌HW�C�rY�Z�|�X:0���M�:�"Ա�����R�h�x[�_&��|%L^�F�S� pU`�2BȜ��S��#��x?��C`��)A��%��|�N:�H�{]ݖǷ���v�I�N���<2?��O��P?i��R֗BT��?�+r:��������n-"U���+�*
�#s�_Z���aoL}*:��:������L�d�َx����*GdĘ���?�,��|�ԢR ��P���FE�qS��� ��#z��|��]_�	F߂� �l0+#��1�+�g0�V?��8�U:>Âi�ؓ�E����^�W�^�aP�V������+zGw�
�:��e�L�Z4�U�I5t�TuG4Xt�u��O�TMx�mҨx�Q�74��H.�`3��H��	����e�5�z�3�G	�?�m�!,��4�q6����7�K���/܊-9��n�r����'��k@C%����d��F���6Kc_U�n�]V)xh���S�O�  ����C$E�O�֥��yԋ�0� �Ghު�����_s���wϭ�,�PS3��0�')2d��1�w��_��~�OIw���JYqH���- }l)���70zt-
���!��.��j��G��=��=�Uwa����%}����;@-��M@���+�.;�F��B���	��d��ҭx\n=�l�`�r�K�#Z��������8�#�QԄQ�2����9'���߇ ��X��bBc���t+�hc�C��̋ zo��fbH�����`A;in�txV"���>Y��Z�?�p�S<�Rg�x<��H�?�Qz����yð�6ɞˆG���[�Ѯg��T�6B���G����ZEM����ȥ��:NJk��FC2�H�*p��'��O��
��&/ć�HS��Q&����1r�������f��obȡ��B"�^(�_'e��Vg��s����+��N#�����	S
DQ�'��fbn�6��H�(���2��[�hm���m6�S�Ņ�sk@��醴3g���2̂�}r��)�E|��\�}1{3�zH��������<���7�tD)����#J���Z���dW~D)���]�Od�yߞ�����.*�Y{0\g�W��H��Q��]��롋��<�����ȣ21kN� ��(��yRG�Tl$:�=��!f�+|����q�t��	�DXT�����V��!��ϔ/w���fI�V���:��CX�$a��;�_���a�
>��V�?����:	9���Z�t�mC���g��ŞA��u��n����J��V��QhT�MN�T{Kb����:s@��2,��f�#���r�Ъ�4�6.$=5���ٺ�Ij�~��?|*��]ܭ�$[�ЩBJ�Y�k�6>ZSF�o�=솽�b��2ٛ�U��nم$�p�&�Q��al�g��DJI{Llv4ss)VJ'���Q�CNL��5A�������*Lm�L�~��i��P��w�r;�+m��M%���h���vƜ����6�����wA�$zN��~��z��E���&|���L�A���1�yИ�@��,�?���+ֹ��Vr�׼�0��t��J﵇2��-���o�6fVf�i���^x�l�q�BQ�H�{���b;�|Qz��i٧R�4t�5�;@�+�3���-q$?!I�3c*�4��m��?���7��4	 �J�J�n }�w����]~4���s{wl���qn���܌��Fz�0~]�>�����$\�JZOj�n� ޔ����B��Ym]��c�z�֑ �1�>��s��*���8sa����d�[��i���kPI5�C�n�+R6Gə�lw�ke29a������kB���Zi�"˥_\"oq�s"&�C��;k�Dqc�#�yx�B]PY0O��y�.= H�?���jz�Z�����q���W ���U6�a�ޞ�=�%�,X|Ϙ�)4��zQ� \��6N\���ɠCw�����1S�r��z�!�V�)pD�5�yo��aђ��6��w�\V�	o��)f
v���{f�N}��F7k�{�jPFe��+@����#f�6�������8����Ɣ]~�DM<��|�x��O�Wwp��/������H��h�E��f�]��[���\�qԫ�f;�����¼˭V�@��^�����FR��`r����.g����)�݆A�����}��3aDyء�ĳ��9Z-��RX6�������K��LT28�|`+���|g`���5���9��);�O6�m�Y��B�2!0�k���qQk�B�چ������G�;Zʣ����;]a���J��wRsk���!���҄6m��-᱌�89�i���8?q���)�i���Ł<M�<��ڪ�-5���5�F�=�B����3�ʦ�#sq2�I����f���M�P��B}���j�� =��pK�Z��H�T)d�V��#']$���B.�271��.ti�=Ug���}Bϸ.���lp���a�� rO&-�Ir�ǈ|e��;�����F�xf�Zޤ�<k����,�B�ҒU���ՙ�&$~���vs�yO,�^<&��U�ô���A,&����m;�]�X X����@��N�qHA� �r�*�o��5qƓ�"�t0'b5|pO"<K��y��e��ݢ�=#�`��.t�����?o�8��s��B��4��� �h!�m�H�Ri����
�ą�5'��`�z����O@������Qwa�*%;���](�����D�?A&[u��� ���dh���T���s����>��1oq�/��I���Y@�\q���)�.�>��I�t��&B�e�p:V`�J?�=���٪�Q?�������2t$RO����aL���k}Bqo�VԦ��pn���aW��~+>��n;�;(\*������&�XT��M����D�!�ϫ#�r:�,��b��|�	��L1�������'��v��XI�o�j(u���*tasn�:��%'����F}K2Z��@��ih� p՘�UJn$#ua9U�j��'�	 �*�,$��ז�!���TT;�KS�D�\��*(�*���&8t�X�}��4�[� H$�&=�k��s(��"����)�L�	��>(Lz��o���G����Um#�]��h'$W�"9���Q�+�� F2O��[W���Qޙ��5_�*_�S���Q�׽���K�5^'�ۑhP�W�z^�~I{���$�kۅ(����я�){Ԋ���O-��%r�t>n�AۂC��;t9�`�_�6�
!@���e�`�y�	����+�J�p��^%���ܲeG�A0h��9R���A�l���L��R�oF��+!	�iΟ.6���x���o�-&����օ�	\)�%����L9����~�Ov��YT�^�L�&�a�lH�P�׊F����)0�p���9>X/�� -�7I�����k-�_�h��J."�	O`��C�F���6H^"hgJ�[��ʫ~E�UPV�$&�74���b@�nę�k��U<C�ޖ��:�p&уo)�y?����`�!������3�\lc%�3�@�~��J�kƙߚ���v�C�J��&3�9b1<��3��ȶ����{��Q�@��WI�u ���侽:�=�<~B�rL~͚c햡�$3�HL2m�c�m�5z�'���4�^O�r�Aj���L��� ���7X8�AC�F��ڀ[Z�Zp�X2��D�����������[vƳ>�:<��&#�T�x3,��Sg{�G���$��`|�96|DY��a��5v�7~J$D��i�1�Y�{�ԵX!%)��N�$
ZO����T��c�������ļ=r~�"��Z_���[��O��_��� �����6:�I��4�T	�,�`�*��xVsK~w��*�z��v��o��
��^�΀����{����R���e
�^�uje�����*弆���ʩH�/J(��8~L
�r��x� -�6����x�]�� P�l9=2%�Ie��Zv^�J+��9"�ǽL��du����L�_$E~����y%��z��ۣ�+��?;�]A'C�aM�kR���f?�u$�@�,NUsC�Sn(A�j%X+��W]�q�^]��䉀ʔ��U��.״�U��%$���e��̬�츝��2J04<���G�9�Nȡ[�V�VZxQ)��3E$��\W$:Rr�����qh���~I��Đ���}��96�X*I+D���wM��H^!u��|F3G��A��\_�wa�����|/�i��;a��) �*�YT{2:B�R.��	�I_M�L��q��j%\*�@�B�(J��4e�ÇZ���I�
5��$5f�)B�>t�:Q2��}�ac�g�(��*%��{��}˓(���Yw�0�^c-ܢ�������$�����\w�|����S^h߲��1�`����3��R&GKmj'��g�#�F��K�PK�p�pJGr���qÈ�H&+���릹Z&��j���S�s��:O^�D�l����k���cDoP�R��q`��I��|'+�Y����!hO�Y�g8����(�v��'H}'wt�$�j������q��y�~��آǴ��ǉ3�9s�`����زu�&^�_*!_�1��Mr�����F�Z$H��Jx�O����`P���S���X������ԛQ�ڸb����(��~�Sd������#�EC�d���j��g��1pBx&��c��i�\yr��_�f~>a=y��,�Lw���跹��@s(�O�CB�w��@�_��+X4:^���yR��R/GKイq ��~�F�Shԑ�X��|F�8m�K2�sF)�3 �U�����&��nKi�K�L�PUS�e#��a��Ke����։����O�;���\�h�#b��d~�k����)�L�ꋵ�OY"O��{�p��wS[��w���̗�th{��R���$��$�Q����g����p�g���{�Ը`��sD�[H��8s�c��f�+V��y:��� K�"��Îx�.��� "�pu�Aߊ�̞	ٰ�Y��5��LDGNȀ�]�C��8
!(����Q;��{nVl��_��~���g_����mR�^m%4���D-�t�$ �����������T��+�t�Hm����}��<��rf��jf�fDC��Q.$E~\�.Le�K��
����$p\@����_���!��&��r /�jRw����N{b��"�H�o�;�����_�OP&�!A�lS��^��6
&)c�@���
�F���9��;��p~�I�������^��`��:	l`Bf�mG����2�ւaht�KI�9�mRgZq�,a>��J�?�q�n���q�)�=;鵘C���zi$.J�}W��f�Y��*byǿ0�oY��d�ڜL�g+O���,��2�E���:~�L��ij)���nZ>0��q�(?�S}.G���(���*�i�A���UZ伧x0�Q��um͊��u��G�����.I����2�#�ϟ�#k���������-�E�`a�fT�)i�ay���o�5�$�!9��@�+�O�!Gw͹��5���]a�x,l�����~C�[)�<J�)�K���Ii�=�?cg��Ut��^!kT%���OTggB�\Bt�NsCl �Y�b]R�i��ߚ2�=��Y����H�nxM���va%��QU��Qs�y�
 �x��E�"y;Y�d=�S�W W�e8#�(�J,���>1�/���u#Q�/��^-��MɊy���h�c�'��
�g�l�ֿIS'��� V�Tq J�-�(�0���Rz�}U���]�����Fd=�N#�����T�`����<�e's�*�=���l�>� ���7	� HAP�C��-h����[�`v�fA�}it��0��E���C!���U��3C���4��⶘���f�����c�(���Ll�w�6������6dy(��e����\m97Ip]tY�Zb��_�ٕ���9���r���t��_롈� DqC�j��h�A]����j��	[j+�wӳtp�|�YI;§�f���� |�Wq���`�T;�s��g)�+�W��E,�(@������@5��唑�.&��Ck/>�L/(	� }Vd��/Uw��,J��P�����#{%A�l�������g,����l��مYخ@'d��f�_^��|a��'��{Dހ�]!l1��!�O.
eճ���SMx�&X��l��V�E��v�	����5&^�7��T�?���l�4l�tj6�簭|.��祬����	"g��q��3я��r�N� �������-�t�6�z��rzNs;5����w��0�~���y�Xܨ���������y��y�'!��3UQ.��V�W�K҅m��˪h`^=��9��p*���c�ŝf�rܗ�5� g���np�oD�g&1�kǉ=�f��m�U �v��;1fH�&�ȞD�I�Y�Na��-�ߢ�Jv�Y]�)�0=ne [vg��wǛ?΀G�t/�$f���	2�U,��x�$4������vt��^�����s:�!�υ�CI�D� 4˃�T��O��d���>
ɵa�tJ�8��!
u˕��.���
A��u���	��Gv�4�jz�ߪl���+)H�g�Ξ��S��:ŷd�?��@5��x���i7����P������)��Y�*�q�Eƕ4�Z�9�p;{7}>�0Ǐ�kT���I�n��(q�n����G'٦f���$�5�vW@��G�4ƪR�%�C8�
f��7�P����_�Y����U��
���A���e��Q���G�&�t;�p91D^%fE����n�G�zױ���!ŶԼO�[k��m$pc�t`�Yn��`f��hGx[} 삿^n�D� r���VN���v^O�1j1%8st�;J���1��E��B=o?q_��j��ɦa�-�"7���<����`�����-�) Fk�J�ҵ�݇|�"N��?[��Q5��0�����%��#�ԉ(�փ�L��(}$t�2���1�]�>퐏��L�jѡuhd9���_����2%�E�i.g(�kZ�_���!�a'O(�z���ӘT���Nd�|ED���T��Sx�-�UD����Ϳ]�����^Z�a�`���b�L�MV�P�6�j�̱˾�W{�d]�Ktӡ#�Lz����G����
3t�q2������z�6��s݌��)�nM���Ӟp���`�b�.(��2ό;���aO��bw\�<]�GTY#��Yy���h>.�'jO-�e��ʧb]\C �>��c�bRz�L�9�MХ�^���u0')����|r�P��U����y�L���[E��{��77�z)��7�v�����W�b�+�dz~nE�`��~ �;�{[�Ϥ��,�e�`t��,5��B����]��B����̫5#�6����]d��ߖa`�D���XȒ�ܚF���?-��fVsK�� ^��9���zny��J���ޜ[ҹ�ʟ��kdͬ�d�vLx�2㾯��7l�6�xq��2��r�q�f� 0��\()���q���^�*�mFu_k �e �v��,B1&`�(��W ���O����i�`��m]���Z޶yÒ�t4Bf�ݪWs{џ�[A{�H�#
��F�CR?�9_��|ȏOZ  4�P&�d7�����,��t��
�P.����g�v��������L�}��T�:@���r��L����`F�S��C�Z^�Q���-dp��IB#��1�����Tu"�ʝ�	X��O\�|�p���߶�&�6���n��Iߎ�t�R")Lx���[In�i.ƀ�Б�m�w������hf���wpM����;����<RTJb5ի�.����u�1FU�	ש�[���.�B��p�w�')-E�m��~)8�tYo��� �$��o�����7�k57o5]��
􊞡X7�]լǾx��aB��X�~��e�v�"�9��k\�*'�C ��j����F���V}�޺���E0��i��h g��V�����̧ɽm�dI�Y�O�����}�^�(ia�8�����lVFO�jǧH y�:1L���d6\U2p�p��G����B՞�����G��ؘx�'���������Փ�@���!��Q�㈩�J�G��4i�j!��T=�e5��BY��R�z�li�T�,�H���"*:�MP@-廏��c�D�� ɨ�"������oi�N����(S��YO����0J��C�c���:�����(Y ��8��A�$��L8���R�{'�$�&��>H<���a��e>�Ehw�+Jb3w��^������O�<"���Xyg(���a^l*�<��ԊU��B)?UC_i�^);;4��T��L��P���JY�h40C��7� �眊ՙ�HN
��	vD�>�q'�/�@Ʈ�Q�ߊpH"Do��9�i���a����Ļ9k��pg&s��vXl�;���B�����r �}j�{�	>���	�Z�1KW�U��ФE�zjzK�*a�T�7;TRX	�����?~ʌ�5%rǎS:R���k�o�����Â�7xU�\�ƕ�jrUΪ�����ZS�z��p��z�%�OG���i:����i�Gi�����|м��̤�Ҝsf��'�*=���:ͩM$��x���-`��r��� ��l���3���(Û�)��u���� )�&���>��7j��^���O�9���R��S��<��y��4��x0Ic�S�θ�)�r�Tsע�]���(�U�ڈ��,~�=Ogéש�g�J�B�-%B�&�[}	������f����@��ӹ��N[:-�F�4�m-��p /j?ia7� ��T�73+�u�m��x�\���H�S˪�.�_U��O�3X_2���_��i�[����Y��S E�+ZB?��Ξ�Mm������C&=	�^������-�PK�j����@nb�0�pi����m�O�cyitճ�D���R�y,�'� _���h1M�8�kq�R�8:TQƳiܢ��z��z�v�+_FH�Im��o��M%��R�U�o����
v*Wk����M�z4{哏��!qʉ�4���)�u2��m_�� 1���<�!6��DSἕB�8���k3�z�#�S����O����7$�ܬ䦘��7$R�"��l��V|�t3ᛈ��.�f���]
7�ĝ�������c�B�tC�uyI��R�(6ze��c(���ĉ:v.E�X+
H��zo���[�N�����6��������h�w���O����ܥ60ހP>_�a��`׹se2{|Kn����Y7B�5Al�
c:��6��=1�ah�N�8>g4�`��h>Y�/�0t�EB�8W>��0Umj�.��HׂLz+C�8�WB�&I��F�R�@d��H���<g�Z5�b27Շ@��C�.��x�~]�X�!t;E�Y�f�A�vx�
�O�<醊O�s��Q�E�G��Mp!����8x�:�8��ٲ~��R!��2���(38�p:NDtcrä�x��u	L��5�� �o�j��0�J��=�W ODr8�(c~�5ں]�/��C��`����E��Ʌ�r�.eui7�q��O{u���D���Ė�o��v�h�*d�mtݣ�]UG0	��fypa�O�j�4-^��-Q:�ʷ�f ��a��(��m�h��96c�* =���	��D_�!����$����=�c���CVC�^�;�����ot��Gw�F�8��>��l2�lL1�.��ғ�)5�8`���"$A����/q\��@AC�Dm��t����,��炓aÜ&A�+jAQ�F �9;����PZ���+Y[���� Z�g� ��؄���_Y�v� }FV{�hx��.� ��
a�:�I	�r ����A��	 �_�&,��I���5�����6��9鱯*��rR�����W��mϟB��S��xM���Iei�;��X3�:���Y���5&����8��]O	���}WA݂Ҿ�n5�ɝ�g���Gso��%B����`ph*��!ߴF���� )� ��5/Jo�4�����3�u���;�l�{�6��|�`:�����BA�0[�u���{g���ѽ��OeeR8��S�#|�	)���ķ}>ȞQ,��>�_������GWǘ,���^�V�K ����l)m��_�Ȭ g���+ø���ɤo)���ss�6�({�t|��+
Ua�g�i�(.\7d��
ݕ��ߧX��F4��LJ
)ƒ-�����h�Ӫ�%A��[�� L�D��������l���qt
�m�xHW�۽�>v̨Lk�V���%���m�8�#	�>��2��܇q[�,����:�8]F�@WS_���p��k<�+վ
�{i��:�f{{R��\�(��N�3�͕�LD��>	�h�Ӓݮ������ۿ�t���he����Ae��ZG%ډ�m۔�X��A��������hW�X����������� �* ������Ya� �^�0H�q]Y&�^�o���%�m���ʁ"aڀEIoտX~vTa��n1��Cn��كFy�tY��t���2ڪ強��M��_�����"�y����Ɠ��5ޞ��-&�!�!��KLnQ�F|��3��A�K��z,�z�C��� �z�E�U�I��W-�	�'<y,ð�Ml8��*�&����o���)t���,N���[��rc=����{l':__`�L�N�����AL�P$���{�s:65˕�����=�\1�k�s �#���H4�9�����UI����{�^�!6p<�!g�l/��ZSHsD��B��8��Dm�3ih���<�X��Qܶd��.,��7�������?M�7��c?�[���n�R�w!{A2���!�B��4��@��v��FP��F0y��f�h��Þ�TB�1�l�Ԉ��4��S7q�C݉k���U�EWf��hW1��9��Ib��V܁ީ���M���P �}H�u�T^F������������7k �{6t�KC�xɶ��&<�|���6����͍�����e٢��lrgN�3�����:W:�:� o����*J�Yy�0Ycm�L�欸��(��B)j,,
9%��I�ۣ����q��O���^Z�.���̽38{4����{����Pm�	��S%Mn����;(�gY
�\Y��9).�.�ۄ�^6�
v�|���[�T��杻9�㥥+&w�ba�	-��<�K�����Z�c�n��is�8p�Lk���4r�4�P��.%@�Nu��	OÂ��x�W�a��ɉ�W$�����5!�G)V���?#A��~~���l78�P%C�D�����/4?>��:.����T���_���C��|��B5l���9�,kC��7�-B��K3��Z�x'\�|�'UuA�M����x�>�,��G��b��f����>�9�4��LF6�(�YP0r��#��d��+��=>�'�+�3�ޅZ�J�}��5i����gf6ф��#/&�,.�ToGlTB�����.��"��Ȼ�f�<�,M$���C�<���z'�Qq�ʬ2V�2~��˩�CB�;w����� S�� 7*�~��g��#4�n�[L�e�;N�P��'�@I�I�M�o�W��A|��[��>k�֦R	�������Q�@@5�0�k����g�31���̱�t��ݫ�D�b eb�����c�h�n�׶Z�2����=V3p�U����i����IL�I��t�X�R[�XG���V�����1��A�M�*��i6B�8�� N��kpirY��
u4�`��h��W�}R�%`Uxk>4�K�ۈ�73��� k���Z��;�~���q%��Ug%�j��3����SΔA��d�[��n��>����i�,����2�Ǧ?8+��*� r�i(9�@-2:�"F}��'�=�n�"ym���T�z�t6"W(�_�I�s�Y44 ��k6��)��ᙺ�.+'�$'^����d��'T���f[2�;�w%,�h���[%�5��HmQ���y����^�>�l�Ja�+��-$ ����W<D�/W�X����]��z�+��,�=d�?/�(�[�|��-�f�,d,]��\��5P�g6{6#�'��t��$s �i�
��y)G G��,*����C^Dye�ZP9��$&9ӵ<o&(<�����3�9
����U�����Kn�m��Mk����x��9cZ��ksceĹȻIq�e5���=�5�LE*�����gGG9P�� �����;��8�c�]��s�o����hX.C1xl.i�p�x?=v��^Z<�᪻����$~�	1��\ъ⩔��Zw#X��=��R�b���ѻ���GH������h��i�aX�;6�^7���]/Byb�hJ��d�_����`NY��1�l��B?���̒�zӺ#���P�����o|�y�ZO�[t���N�>^�'�`]ȿ���[�|���n�e$5(����P&��n��l0����F�����/'� ��%�GQ����(�F��Ys���4o9f�����*�\tT�6�{t�Zݩ���SvH�I�	u�P�(��?b2�E�i���%��+Ѡ68+�vD$��	�uS+��r�I�2w06N�� �3�E:V�Ԙ���C,�g�Y� W_<��^�,���6�
X&릂�5b��K�H���.�a�G�9���j$d�,��KY���$j�z0�s�����Ŭ'zF����pś}��u*茢&Ǖ2bč�#·�������~���ș���w"o�Wc} q;8��b� Yʰ�3c�1fA��Rp�9��/كXQ�}^w��WO�=���U����=^$G|֙D��h�gNZ�3��L0CPz[8���6{NN�io��<af��@�	2o�n�>����^.��A���'�{$�] M��N��60��E��U�m�en�r!�e�e[�1,�>T3�T��(����YĂ�l#g������������_�R�r`6��fМ$ay���ʵBuȰ���il��C}��V�~S>l�&�mR�(��M��k�S�,r������)7����?�la2�Ir���Do�:Z�:p�*�_�o(\j�T���J����̾�2�p��b����� �"m�Ȕ�o�}j�6�����.�U���\7�zJo���(߮l��o�M�R;���R[ō�͖��s�æU ���3c��p�XD��8ބ}��`�S�u�'/�͎9*�WP��eLy+n��D�I�~�I]��Lyԋ�|!%Ԧ-�W7!�ՙN:,��$*��	��Df]
��:��ˢ���I-���þC����摣� ��b5O�k:$��!��@�]�k61%��$�5�c��,�4鋽�)l@3yl�h����+Y��� B��Qυ얆����`�����?��F���oj��z':h��5w_'%�צXǔ���j���}&֖�t���{t� -��ؿH����ϑ� ,m���O�����c�$�O?�P���3K��� *t�J�:%~��D�*��ɩq��`���XON_����fuE21�ƒד>8�KC]���8�������tp����y���f��~bP������3aE�k�NDΆ�{�X�<-��O���b:>�QaL��|o�}���+�Y�È�3#cOy�zo��*��rrG�i���(�qNH�?<!�� <�>cc���cu:�}�AV}�s�u)q	��[��z�*���å�����΋������S2�F^ƣ8����"PA�5�E)���xp������.�rYC��L����r8u~�:��Q^�I�,Ө�KL#[7�n�'l�7�a>�lU�ŏM�C��p��'���$k�;��e����cf����2�ɱ�J�f�o���[��"�׫�mL�B.@��$A�SPk\T�8�?��;�`�hz��x+�86��~��g2')�w�y	U��X`�r������c���qO_�U�mh�E�<#�젂-!J�������aS�e-��0���TԕJ��?����%EвI����s��O .|ɬ��Yx٪��j �T�=���ܝ�x�0��>ƶ�{�Q�����zv����o�L��K�>��9�
R�{�[%k��5�-��8�ɥ��>���riX�`g�ڞ�(N����7ٞ�ho)8?�s#S��wd�Y��o0Z
7��h���qZ��X:�mN��}J���l�n�q�Q����]�ΛFѧU*����&.��-:!�|(:�2mR�ME����� ���Z;EA�cq�U��mȩGx�j�e�D�$Z�"U<��-6����1�v��$�;8�H\���D�u�M����ֵP�@��E |����dӳ��=��}S$,�˖��j�t�Guf~���;^��\�����zg��R�E;�W Ѷ�N�sV�� �������NǿH��B>��6�"�՗9 zb8�Bj�)f�Fdvc���==t�B�t���?�u%n��6t�=.H�>�k��a��^��~�27�a�����q�7)��5iO�R�,FD ���m���i��
��j)�̭��v��4`�Hsق�\��R���.|Kƽh�NXG+9���-���~���h��"�
���q��r芒�e�r8wȅ���2��ܝ����rfT�5��E�q�smI�$�AEK(�i�<�ӏ�%�I�
7T�U4$f��v��A��8Z��(���V�y3���QK�
aDM�s��~���˺���� W��k�נb	i�-��i35��짷�<=L�����W������3n�+F��.�@R�X��a��E�\���o�<�� QwĤ��i�z�Q��ue}�k�V���7q�����З��V�rA	� �;.Y��"��V�2� V�5� ��Y��zaz
iDb�A��ds^���>>N��t۬� �6�]��&��xQ�?�?[�|��q7�'�G��3P�ܩvRx�����o���5cK,`J�+:a9Fu
xM?P:P!��x��M���
{�e��LFk$�f��|����N�D�4���v��#�6���.(��������gB������;1��	_"A-��]38g4���-"¼l����y�%���K���G/C5�U�x �7�_��m����d0��Fu�3�3ha�%��Q.��k�9�R�Ŝ�������؁��SɆ�q�&�q������b�>pG���;�x$8�?��	&��/�֫�"�z�4�r�}���H��a:$Tf�G���h�M ��N�͹$�sxݗ���0U)ˀq���^s'gDH�g �c����$����٥w��mk~:c��ϴ�7�ܝ�z��* ��(M\������$���PB ׊L�� D̤�{`��.<�ʥ�F����:=�K���Vp�&pP�_��D;$PA�8s+
�.���	��R&�=L&:Fvx�#�m��p-K��	j#j���r���]o_����p{m�U�RPlix3�$�CE�<^ػo���k+&��SB�&�P�Z�A-:kĊ��B.��u+��G��S�)����{�t��z���#:�B����.��΅ ����F ؗm�#��s�토�Y�Qo�D!��Y·�e�dh�4�R!��m�ԩe���n��H�
��u�|�0*��P�<ΐ���POT����50$9��-��9��՜��5@6SgK�N�aG�ݹު���ݼSL�5#�l��ec�(-�#@	R� ��d`��l�y�,i~�3���[�=D�K�ȠI��tz�[�	_��`���ۘ�idub-uT���F���9�e	�$�s*S�b�)�\�Y��Z��L�'p��?��ӄl6�/&ґ�L=�m�ׅ��@KLb��[���v��}S��	��Ҙ�Lån�Y� ���0z���2�]��"�_�I(���������sx]�7})�n�n��}2���x��G}��l�ȕn:8W�_��{)��~��xrf;�G�X<$WU@�X�d3�[r��~�
��?0��T��ɳ�&%`ƳŢrq��#�A�^z�J�]�R�Q��:��i���Klk��L�ǔ�_�_*5��u�!-�DT��VC�T��k`���m�9�����,1׮�~V4F�U�&n���3W���/�DA8<r�K� ]�����9�E�c����##l\�c/�=#0��G*'�^��-`H��p����Ȑ�M��ϋ��hn�����/.˼�z`���U>c�Ii�ټ�$o�r H�	�q"Y���1��	�l�+��#���T��Ok��ǿ��[��f!{J��u�:�v�q/֖����o�$~1�piR� �:�m�܏����!;p�d�uI�)�R�6B��:u��-��W9�V�S���*vw��4�#rdSXW���m1Ռ6���f<���#�Ih�3Ձ���l��ʠ�l	��I��1��@W�� ����_�\&���7�jT���� ���܎�S~��뼧��}�0
�G{Z�����h�x6�nz��-ڹXg�!�bWb�=��L.9��`���(��x��r|:0W�F�-��W�ԭ��h�e׉�F���<�<��J�HǕ��&7DP���C�):�x	Lc�*ȁ����$&,�v��Y�u.]6"�|&;L�L�f�
�Wt?@.i�$�@,�G T��{c��1����S���b�5^ �z @u�	<�_�c�� ��l~>*C�N�`���i f3pz��a��u�zA�7�U��79��@З��;�i���'G��3���5�n4�a��	�a���V�<�}�U�(�J/D��D�U���n�Y����J����*M��M� \��l,��
�:��;��Ò��nE��qw�-h��.NI��A��ʅ�-W�Vo�ե��ػ�՚�L��$Jv���:I��0�h���`ۃ=)ic���z�q}�!t\���V7�[�ގ��_��Pi��-�??A� 'W�/�H�ZV�4���j���(���(�{�q����a"��I��|��4M��~}�ٙ�X�P/$r-[+���M@d�����
���� ��Z)�p=��M�ǧ�i�<f��}�3(��-fQ��#����<�IƬ�4��C)�xV��u���٢?z}nA��;4	�3�����Qh���)��^#�f��ES���%F��֞�we�^
T6�J �2 ��c�Ax�����9%ԑ��?�r�O���kh�� e�E!a��Y������bh�RN�LO�=�6�&�M��~I�縊�g����N�f�e��-��Tcs��(E
��W��;(a���a8k�&�`��x��$��ߞ..�۳q�1ē���]�9��ύ�\l���-:cpw��u6�Vt����p�`˛ܣ�e�p����s��P����`������ʹL���wH:��
nbf�uT�z#)����Jn/X�Rx_
Lփ-��\������us�7�!x��r�G�����}�;��)I����Cx����QUB�}�@�;2~���f�1�_DL��}�#w�Ş����J��u���t���j������V!�����-��z]�?4F}Yn��adk���P���;�"�����B�p`~O����wg��1�|��A�"3��3�DYi�)���D�t*�A�6���>��YrY-*�,�0z3�'��88S�	y���3����6��.�W8�&޳�\����v�ϕl��w:�P���Ի����T�/B�=%�2��(�4údr�qq��m�5e@����%7[�sz�P4�J��D�>C9�M����;l�B�cj� h���Eb�%4k�H�/͕�JR���%�|�X9+*��'e�ܤ��KC���9t���&^&q�׀�Sq@t���v2����T&���\|H�4������m�4�q��j�a��\�hN���.���ea��`nPKz��G�!��!	*%y�I�Ԅ�@ϙO%k��Y�M�9�I|o-��"81�����w���{��լ�O"�h��U䛌q&U�X���ԥ�$&�^�X{�}-�����i�}\{�ZU
�%y)dS�V�Z��M���v˧��t���iB�\���E7�-��Ƕ&���5�9�VCB�w���y�C�>�**L��W��72��r_�+��|~�z����a{���5ںx\)� "���-z�A��qlK;�U->,�����SW�D����~.��\_�t΃�b�1���lԣD�\��r&�a��_����Q��|R{Cq���S
��=�3h^TLr����<���S!��<B��h>�;��Gf�-⸻��E���=?��F�1U8��z�{��؜l��f��I��-������8�ъS[�k'WdY (�M�&�Ԉ|�k�'�e��c�4Y��_5�MWP�8[+��M����chCVU.���8��$B?������ݦ^4����f0d�FJ��`o=�����+��E��#{+K���q�����"�	�����2��	vU>���/m��k���}��g��\�E��B_�# 0@��|8�S ����f���u�anm����RW3� ���z.�c'�ݱ��m��B�5.Wb�Lso����V"���we�;�40��(F,����a�U�h'n��<;���kO%q��+�3_�j$i8��h��\��p�n��#%��& d2�r-<�0U�R8���F����"[?���d�I>y�cY������F�
��2���6ڣ�{��,g�튴Q�=�r*��?�9��ko��-��p%�:m�Qc��6Wd=� )n��.�v	��%<�0��ePQ*�M��J֭1����?kt��!c�� E�
t��$�g��/��~�Wg=�\7�4ȂE�Rh��&Z��q��43/���_�׉_�/��
��m� �(����Ĵ�P:�:l�p��֚�2&m��s��U[���E�P���YVe����;�R�(��uGS�in}��͸�z������A��K`An�!\��<h:ɬIpu�g�nU�2�@�:o�-�v��eu��dӡ�1�����	���Z$�]n��z���>�6>����%C����Y`�k�/4,͉���h�y�⽋pҝ����i��%�}�2���v��kRq�p��g���
��5|���$�|�2s�խ����u�m�d@�9[�"D�׀u�{��F�Q����.v �Y��ܤ�#~��j����M���I�MZ`�в�%K�U:�`k�l�����aX�v�C1�ց�jy���\:����e�������k-a�@�����`�Či�	5{�(Ӥ�I�'�q<�2͒Q;���>h�.V(t_j�a�#�z��a*0�eXP�* ��*>mϘl�T�BO�,5/��L��%Y>p7���Xo�Oa;iT;A'E��2�S,͘��>�]���f�����]N�g��ܓ�9PkV�iRϘъmi�[���IC�� �W��t��;*1f��O�F:���� �:M�w֎����В�)ʕb����@�c=�+*�re@�V�g�c�g7�mD�{;�k4��W���<�h�ſ�����.�N"��9G�K���0r�DЋ��?C�d���fe嵺��֤EZW�}���i�4��^c^"Jr`_q�鸲6�EI��>��r���ȑ�g�'�j���Qa�I��i�b�ԅ�l���=)�p��"�}ڢj�?�G"�$e-��6�A �t:_xt��q���f�gq.��;�]�E�4Lv�{���L�9��
-֨�G�`%b���Q�'��a:�K�O��s�AXS��?�&����Φ/Q[��w��u	ȭ~����Ie)�+��zr��ϋE��c{��Tߣz�E�<tA���O�r�HTlߋ�T�Bמ�Ķj�����H�w m���U�~�;�1OȊй�j�e�n8[�:�sy����'RL�-����N�N"-�F�tk�������L���φ��R���w���q��R���q9֮V�$޸�hj���<����ƶ���+$/O��`a5�SA�[rR��-�s�8����]�&4ZksW0NƘ&_�12���Y�3�TVk}�ʏ�R����
��Lނ���9^#NM!6^�6������׫f���B�h��K���� ,s����Y�)��{ Z�>K�F�AR��͝�^'"/�'�"��o�F��$m�MG��X
.�ϖ�A!�m#��8�Q(-_��:��0�����,�����y<�J��b�K���P]���~��@|�Øs��t=�僶��BK��,��ܥOI�1� `�X,����ȯ��S�����f��?��dg
�U�#:$�ʥy�
a=��n��\΂�'���u�ʈ	��Z�Ǫ�:u�&>4zL��e���cfυ�88Ь��ϫ}3��i�h�����[� {i �#m�5V!�٧��y��Yrsbi�zc����9�M�K�ϰ��	\É��Se����h�=7'S^[D^�-&J̈�_d�^Y�Z\_[�0T��˿��7��_O��Θ5l�!g���`nЃv�o��ʻ5-�E��~&b^��nb�i%��F*|�j��>���)z�U��_E�n>�)U�ץP�-���G;L�ӊC5�x���ث�X	��(�� ��p�:O3���/p��Ì�Id
T�?�+�R�$6}8,u��44���������0y��hRf��(��/*3N򊦵+�p�g���,�(�%�y�������Rڑ�<�A�&{C�XO�t�:h�%�
:��ʢ���W�����$
����*g@�4��{�|�խ1��c8�* o�/
��JO�s
O0���a�ih(W*r�zHh(� K���4�v�J"G���1���Ħ.���r��Nb�`fA"H"�+SE���M���.��Ua 3��5*�����\�@ܣ�fΓ@�*?�Ʊ��iŶdwI�aQ�C7�,�x���S%�N3�!��CyJ!\P�y�!�������C�/����a|ޛ��I��:�l)���Y����cQ����6�Qi��>�ƃ����U�F��������G�g�6�B5ϩ�*Ba%�k`�R�h�c53�;�Ffb������^�a��t[�"x�=q�#�
{�O����8q[�N����*��&J�H1�+���/�۩�;6.^�;(k�ۻ��X�ˡ��,��\�wc[B�<��b<��7C�0�X���'�7��耧�t�o|&�����'}�p,SK8b8�q���Ên�S���+{�F���#�MA5�6QJ�|a�dr����K������Z��;/�5���I� m���F�B$"���gޯ�&�w�fB5\��,�]#��Z!C��To<+7־��@>�
�2|�=фW]�8�|F�Nyy�C��@��-��$G�2���s��qh $RzܻR�q
	��^�Y+�����V�A,P���:��u����+�M�J�EՋ�3㭹5�{��#b��$T���_/!�z*(RW6�×�	|0�f��.�O�fDEC.��\kU��P���U�; �S���JC�?��J�2J{�C˒����u�Dj&�.��i\1�&M	Yn5+ɋ0+��1��O��oX�Z�.nJT�X ����Oن�8;9�6��3��/�a�GK�<Ễ��Ed֜;:��������9_� �cU��i�9:U�W�2Xyk!dm��Z�ew�K���-��M*�EvaGL�C_:5pk��m�i�`.�Q^U�����8=���~��%FM��m!��5�����W��S��N��m�b-�/����m�G��VO�37@ ���p*��d!�Q�_\c��L��-���Ҭ�����	~�M������W���b���O��y�-x!A��%�_��nh����h��M!�;r���^��v��M�UT��O�����t�#���̙[�ǵXW/�8Mb�z|kś��@>TSuV�ԩP��w{�g�ux�'ؤ�g�V�ݽ�q'f�Y�Q5��]Ѩ�,u��ә8�@\Z����^��q�CF��2,����v��u��/��
_��_��:��zH�������ߨ�)��䍇6���u�vu��f���6�iϸ�|ӕN��@M5Hy1��`Zkz�S<�Owz5o�W�_N�#m�D�f����t�Pã�Z����-Ld��Md��q�������3�B0�YҨf*uG���7��)���g���_�f%�=�\�G�S�d(Tn� �sb2s!��M
�r5;vۭ�QBټmF6,W�k����$��S�Kă�_7��K-r�Dt$q��LE�/0 ��4^"��mh�$�5�y�U��.��#���X� �D��t�F��k.2�7좪����ճR�{�b&�^��i�����x��^�Sٔ9`v��ۛ��u�D���8�$!u;����M��
�m��jU�ɛ���u��zn�V�?r�����#�vA�	�g�\c�zCٝ��-���{����]���ߴ�e4J�mO���=��q��U�q�<Rw�;l���S��8.�U�E�@D�Q�M���@8w�Y��a�����ʌi5��,�������U=����vb0FIbF!�/,�&N(�F��^� pZٜ����`�rn/{^i�D��΄+��N�|A��!�9ß�,tpóK[�س��('�:ʴBSf>�TdD���\r���ݴb����E$�֩���7���2�op0���nF��w�`e��a�H#}��cr�^�´��p���h��X67�Jq�IZ6Q��$��#�e_�f�����$�(�>�*̕c8�s�)�lٶ+!�&X���?�Ø�2DOn��x|�P��dF�r���c~d����Ԩ������C�3s�٤G�L��`�;G�-!.���6�}`C}���v9DԂ��8�m��_?gC��1�#�^+Z䞵�m"t���,�����㵘�kfG���ե���"�`�G[B'�D���`�f-+	�!��/�ZE.mꫭ�}�C�qt6����ٙF�I�.��3�¬]��w���f�"q����
g�M�$n�w]J��'�Vc)I�K�U�XK~`9��W��Ȩ�H/	A�Mtd\��{�C��΅�M�R�/V6g*,Є�x���镊Z��vl�U�^�N�|�}�&�����|A;%wɜN�$8��?.�p�gy�5(��M��ٟ�qy������+@��?TFÒ�!kV�q	��d���Z��Hk���ם	���l�?G��f�
�[��_�z�_���Ⱥ�s���+�����&�� ����
f	x�Ʀ�%d�����J�AP�8����|\�K���M)�z@*�FBI8x3egɊ���o�辮uK��H�@����ު�f���,� m���m�-���8�[���v�Qo��x�si�h>��#h�DNo�b:�v<�5m���
+T����~� �����;'`�����k�E�vm9`�0?�~R��1�+ɶBjm��#���У����nu��'��]�R����.[�a�UW�vY�RL�T�SY�*�AӒ&k�	��,�s-��J&E��7�?��t8RkÈ�8�/L|�8 h#���7�Fm�a�I��-�B~�����d�,Ƀg�����r�r���r�a{u��`���'y1��8��+)�ه�(-�}���C�m����stv��px-�b޳y1$�}]~	�/϶&��2>C��$jX����=n��5�Q����?o=�B���U���
 �"s�[ط���J1�&*>����0����$�7~"�}7�1����s��b���17.�����K#ߣn���T���S�����A`scY����nu�P~�`O�YoY�"�%�3�I��g�`w�-�ϹY]���.\Zhy��e֯p�6��07�<+�ߑ�ݟ�@�w���v-�gl�X?MYvO��T�c�؝Z�'P�ĝ�����c/b��LҨ�{�C�:���8;X�㥜������ҎJeZfvt`�g��*�D�t��M�C
+���ݢ0�q����q�z(�j��r�:w�^`�/l$��W�=���I���kF�m5]
 mm�K����"�>`H�_�$��'��/��!^vn�Q�x��B���I���ј=�a��??�:b^�eU �aj�-���.Y,r2���]�rkQ�	~�dv��<?0;Γ
�r	z �Ԁ��ck�ʸ��X��0�6����_���Ko�]��A�!43J����iS%�5��j�FF�����P�i*h�>م�o� `x���7���T�8@�#����o��}��&��Q�q��$�p��l=\JBt���ڍ"�
#ܢlq�0��p�ʄ4�"�(`�������='���py�e��tBzc��Z��KGnY|-)���AލiZ���^F�x�ũ;���z�z}�n��y~�(���򴽭P]ދ'���U��p��ú ���4M����zF�

��s�����"n̪�[Ey8�]eWW�3s-��Op���c���Fy��:��ek�m�&�Y���,��z���"���ض<�G�\^�Zv`&����g�f�����:\��}�1��fwPmjK�VM��B�s�l��t)��gk�Ӭ5�ԛS�;����O#�CfDs���g��D� x���C�nH$�}��Mcpd�[���Kb�ѥ��TW�ܺ�>?��*l/�W��1�eB�m�ކ,\�#�siS��%��DmtW_�>��k&��g&�!�t`�����Q��N6�H��H�<����?�》'�d�z{�N�R�\0[��w� <v�9�ǌ��6�����Z���H!%����\G�ոs�K6b���@��!�ϴ��&�\+_��˨ld����K^�8�Ю|�Dn�vU}�$���}���&�:�����;��-/w��-��g���2`3�,V���h�P,HPqcӚ�	�m�����[ VYx2_�r2�&��4Y#�Ul:(8WO�����	��n�-<6�< q��ˑ5׿O�	~��4���hu���ꄏ�7��ɱ�8;]�=�':E�7	z�ty�����9�s�t�@�S^��«�
�q.�toǞ>'��Z����nSi<�$���I��y��a�Q	&��e�|' �a�����|~O4@א��c\!�^x��5e%����Ð���z}�]~�4�"�����s5��W--��Bm�O+.��h��a\CR�B���'�S��4��
���|��{GJ���=������U�}q�l}Lƽ|�6x�*[ n�iq,Ϫ+����ɔ�����m7`�ǲ@��l#Z�,���!��&��d����qo�}K�`]y}
<��B_z�p%���k����bT�C�5�p�M�B8��3\���=�� ��O�˯.ϨqM�{šr�[�:����Ǣ�����v�*я!��W�nC��F7ŵ('�X��/
P��K�����!�rP[h��EU��-��T9$�A�^��
|4C�h����y�e8�5�We�'Ə���E� g����T�������t`G8�I4���R."OؓQi�c���2�فd�Q�6-ʢM`�k�K Hg_� 8%�Sy}�P�]�?a���-J�A���::	U#���a�Z�B
ew����d4���ǭQ>Rr5��mT�V�Ct~3S��Ci���'����\�L	�Q�b��� 1>ȧլ��&�R�y�һ�_=�3�N-��^�쬩�I��E�75R9���ʫ�QvOh0N*A�ѶY8��ps���Z�<:���\z�
�=�́��N	y[�.�˱�1�4ZQ�q���>�Vr�"�]��l0���N�i\e�q�!JT��+�L��p�ch��&9|���wd����$g�>�w�����Łc�tK���iit��!-�|��3j�-��;zb>.)i���6:�J�|-�$����G�
���d�>W�����S�T/rߕğ5q�`��T�5��S����ב�L&�3��[21<�T#8T@�aw�.�]� ���ʲU� h��|r~�]�|+��,��c����:?��?u5f@�6�q�>R}+�I���KT!��w4+�e.��hV�/#���>0e��D�=���l��?���N(������č��jJd��?�G�I��^�΋1֠�
���#�L��Q��PL
�]�1��e�X(���ܿ;�^h���/�0��y`��p�G)J ?�1�8�h:+�����Z{刖�^a�i���3�A9?&��9����'�β�<���-w�;�6v���n�be����.��@j_�#�!����O�0�����X��d2I����L������
�KLu�)k��Shh�R뛿B����p���:���ض��V�,M\�I��x���	v����<�^ܛ�^5�ʊ�?�:�;¢!�(;���*��6��ig���N[�#o�{�C�p��t|�m�aL9��sBvAwN�v�`d��y3u=�F���1�\ ŷ��r�y.s�����V���ؿB?�Zd�5� )���a|�A��\�tP�U3Vڼ����.�����f��-4�i���(��gu ;?���G�>Y�W�O�F������G�ު���IC�����]���{M����WW�t� �nI���xq�@ltp@�ɛ��3�҄�ѵK���k��`α�]�^(%v ���?}�A�.K�t�Y�C�!��(s�cf�y���0+(��� 	L��M}t�b+�,�i/(�?_�#Y2t��9�v��D<����h�H���Kl9�}R���ܓ���~�j�^|�_�;���k�*��8��rԭY툡n�8k����a��-0Eג�5�(�6<�Ttלګ�&��Q��1:�;��>V`�` ̈́OD��-����|%�l
'��iU((�R)x�O��nE� "i�$�0� X���&rݕ�m�2}�H6�p$�mȑ�9�Ϙ�΃T��Q��֡�i����'�8���Xi46:��@FG��g 
0��x��)��2��B�
���1q��N�ߕ���M���a���2�K��@����͆�y�y�%�u�z`�h-�
ɉ��G�
�+ל�
� S�/�3i߯xh�CT'��Ek�/K�c)�$�i]_���T'��7�f�כ���b����7��"n�dxpW����hN�G��C���(�M��d�$:ƷE)N=����93���gޖ� +��J��)G	R��"�J��>ʓ/�=K��^��ўg|��I/�Jpۗ,.�8U8B��1���u|Q���YLҝJs��0e°L��C:8��g��(���L���@Y�+� ���L��hT�j��hp^ubA�vM�c�|��*�\Ő�J����4��}1A����8��Щk�V��bSD�
�e�Κ7��
���!�'�g ��n�w)]���2���lVh,F��vrE<�"��#b.��i5�e����VΎѣ��l�1Rbf�oE�a�>�OC@�m�����m�Oc+7C�V)�(�{*�i)��+�h�Ѡ6����B	wQ�~)��Y7Rb���9�ݤ�$�?��֜3d��rl�֚a-���b��K2�S֑lr��l]*���m9�i����)Ot��՚>�ȋ�@J���6���:�.5G1ܴ�L֕��E�LXp�RI���#�3Tכ����j�5Ǔ�&�ĹX���yL]h���PvUB*g��10�H�k{�����s����3���.��,��_�.�D����D[	?Y���"i���y���ѡEdC4ة\!p�zFHr0�0�?�` �^�'i����v��V��P�o��9
�6"mw��?�a�0� �l��Rq'N��_О���E"_q��ۇI��]W#{[���i8��Q	Z >�e�3��Z������/.��\��g˼z�c�<EZ)�U�ա��ԽE��o9P���� �?��(�`$��;�A# ��_�HA>��%�s��f̦�b����t<�=�;fMm���%.�{���:J*s2� Cb?���`<���5�J�'�#�,ͱ�O�����)�4���=����sK{��P���*~�����9^,J���fe�!|����HӶ��p�2�kǶĚ��/H���x^� ,�R�m,( V�n����b[����}�[�,~���H,�6�^W6f�۔����*]�EA՟;>�!1yv��-M�8ky6��M��F��2��wǦ����i��ྦ�v:����{��02�_���*\l��Q)�s����� ,��tp�3�&P������K�s�����I�4W�#T��Dàp�̏HEl�ٵr0?���*BZ��#�!���$c���I��<�o�W�ݮ��Sg�|���C
^𾼥J`#�<�t�<�`�c�ӯz�]5 ��?�զ�\��ߣ�W��"�/�^Vz.������2�F�&�I�Te�R#�԰�����Z�2��c��]_�1��k�st�z���8�>[w��rX��ӊ�?�Nc�l��C���k�7�<F����X��j�hY��L52U��a	 ?�_]L4Y'��`�Z��䂅�|`^0d���/����>��`&�b��U�p�	�½xh�3�"��|?˰��ծ��8q�;k�Q %�5�W��b��77�Ly�R[h�TU���m9F�ܡ�Ө��o���o<F�["ڍk�]�lN�	�T6]C��%��&E� �z(�+8�5[��Y�HN���!�Q駑ӯ+�rcs����a:G90}{t5d�j\�P�o�Vi�d�8������c̮����3�x"��'�q��!����o����-����t��O��Urk�8��x�S(B�H�N����"+'Tu�7H)�����ge=X��}
�9a�[�:��3һ�ܞ���Se�<��F,@�l���m��# ���G���.���u!�N5���E��\��Y�TM|y�O,D��@�S�s����� 4�4�m���)�YK^�A���$�� L����ڮ_0A�V<�ܲCG��,�Wg�K0u��GY��$�즊!�AH���x#�r<2ӫr_e"Әmq7�)�.�9N,��~�� #�5���tu"=3!I�L��OP�k��~���O�^\��V��T4�u����o���A�Y֡�V+F��W��HiR���\��PxI��=�fN^XE��[��Ϻ�N{�w�z�!�ܦ���>�9�~ɶ���9��AC�N���7����:��ι���ݧ{]��v)�\���=�n���AG���B���Jҟ���*l.�2z[��9�h�QF�'�T��9����MVz�c���q�����׀�D�����)=�GO��(uh9�?��/qY�kg�d��X�(�m���8�m�E̟p�#�)���@HI]�-�B0n��ׯ$�f�L����wh��~f�}^-�RY�Z������B��p�ʄ��o� �٘���F5��E�qS/H�F�c�N�w���ufLy�K��*_dl���^�*������Ƃ�fq�Ԧ*�VLx{�MH�:_Ƙ���P-z��tW$��d���E4���@�D�86�	O��qpF*^e�@v�zKh�+;n�d��ā�Xo��8��uJD?(���F����]���exh`�E20�/�ߠo���e�=��0���*�G��z�=E����{�SZ��[o�nS����&!��{p�F��>��N���/�dJ^<�1++�$�Bq���
>oLå��,t_@i���Ŏ����i��Gi;�ҋ���j]� o.�U:l^�X���ʹ��3��"G�7bod�ICE�j_�r_�7*�$YOq-�H�wo���v_3�j;�D��0�����*P��lloIp�k���u6tUC}����Be�c6hw	~�r�'��������7^�s���ñ1K�p��"�(I��&M���- ����
��MS�A�X�,B(1���`�q#���/v���4����BS'�.}�˹�{��1NR������̙��;>����]66�����]8�̗�'���'��T�|��hm�H��N'�_#�ln�`�w�X�LG*� ]�j���夸G�8@�N(����-���ck�
P�+�X����8�@7����݅E�_�Z�B��gh 6���!Z<� ��8ֽLAGT�d�|L.��y*7�y�
���J�3d@X�)T�$nِ�v�eL��T</��ط���
roن~�
��y�1����$�&���&��ҧ��b��>Gy�L�옿]���`�aY:�ǐ�@@'��%�����Z4��r�z�2�"��m�`�G���$6�z��o�w�>y�͘�*������.���;5�NY���3`�[[�"��DP��Q���F0�E�f� ���vr�
X�>���bJsi�\�k����H��;?���1a6f���m~�o����`a� Xd�ǯX�p�1G��'k�p���mIf��j�ם͑6r!L����������r��'�8s%$7��E�""��h�)tB4��^����"'�Ȕ@��ڲ$���>3�ݯ(��3����`�Y�qvx~���j�qR/����V`�c������`L��_7H?����a��n}ހq�}��_{]��1�0�{�jtv� g7�%a�vd�hft	���_ф�Z����=�6�>��c.���]B@�B�4��>޸B)�&���^}�H(=��^�-Mj���o5^��?|�¹$V�s!��8�V!y�W1gLI��"M�K��0��$�J�q{�+$pnH�sO����p��GHyMM[y�y��?��b�&�>��ݭ0����I�R�IU��<f\��\#P)�� d�$X�B.�Tf.�F0���hXg�f�.f ҷ�J��wf1�G.tn]I<�`����E�]��d�7k�,	�4��\�a�X~�'ZY���Ny2.��	W7�=��`:��b�+9x�K�-#	����q\��m���
�/�K����EW$��n��=����T�ڑ��⇵�t��V?ڔb�ǫ��|oM�]���{�=b
�V��Eu��k�w��p��J؆�1�@V�Mr��h&m���@�#���w]G-��d���O�]��B�o����� b�V���lq��.�oyLF��C%|/[�SK����yΌQ����jo�K��:�?zz����9'Uf��2��i�5D���H�?��hڜda^	���ghTA
>�G��v��/�H�J��>]�C
�p�8l�\��x,G��KNp��,�Yl���ON��_X�@�{T�����m�'E2&h
�9Q}@���/�H������k<��o�Y��FkV��hߊ�Gjg��:6�)2�2�y���X�iӽtSt�Y��Pz�l�v=7,���=9I�^2IǊ����F��;��h/��W����x5��-�`a����̳0��B�2s�'�-W���þ�d��a�8>]�V^���.^�}�y�n0���R:A�z����o,� ��{Ð�V�-Y��y����6F+�^-�Jܱ�����ʺ�>���o�|v�	�Zȴ�'��ף!zX)�p���d�T�m�3;zko.���l8z,��̉x��x�m����Hw\
���x�����CA���`����0�N#����Ă`��p�R�/{��٦ʑ�c�q���&u��k�V���Ϊ`�E�
�_���=S�i�*��NQ�(�k���]N$o�`^UC8�Ǧ�\�(Y��� L>��ƙזHӅ5�D�ԎD�\.Ȍ؂��=�l1��w�e��vs����7-�6��t>�3��!4���Xаx��!�n?)��a4t�Į��Nd,eD	��� h�9�Q�r���	.����khʼ��zy�N�����T� ���ïX}��x �[��K	k�9�8E^`V��[��U�̐����m"Z���<��}�'*U^]����e�3*�x�MX��j��RƍE��鱉�A�W�3$"ƹMY�ZM�k�'��ߎ���-U�f�`�K<H�j7���Z	� ��^��4���V�2��罝0�}�nL0 x��^Ó�y�¨���q\|u�����ohs���)I��յn�Ns�E�@�L�F�M�������î�2j$>������T3̪C X4�D���Y�8���D�L���>����JA?V�)J�WEDms�	�/�yD���QU�B]���ykG!¿t�G�-�p<���KT�b�\�p�%�ٟiʢo&E��*]hcF��!�T��!�h,A�]��n1`��N��o��N+h��A�(��	[��-os;-/1&�q�]�3� �F�թi!�j��]#���dwO��`�[���)\�;a�^�XlC���34���� E8y^�G����7#L/W�Em]�"���B�.0T`�1f�#W�E�Ճw��p�J�Gy�*y�k��v�慔F2�t0vxw
G�ٽt]��7mI���z:�_cETWl�>��1T]��tF6��y����!J�!�0v*��O!NY�S�r���+n��?�t|h�����l90����0$�.��}��>�l+���:`t@��G�Gv�M�.�{�tU�dj�����Ѧ%5F�v��^;GLջ5�04�<�$��iؿ�8���}�K���,���Y� Q(�4�)�1�~�L��eZ����HRF� ��?h�����<Y���"�QU�ʅ�>Y��]�]�N���P"d���\��c"�!)�z5ԍ�o~�mg�G���@���L!��f��^�H_\����N�5�ܽ#\���<��c��|W'R�����J�+��#|N�z7r6���l���C�2���=��X��|�Z�p{��n�U������+U堢ڵRt6�-c�/�Ε��WnP�{xؗ��\���)Ƞn~o����إ��+����vG)�JWG�����qʈFx�p�bGК ��G&<e���ś��V�cK�×�����4�t���#K��e&RJ�E���<�%%ҼI�Rħ�&���<$��5�hNBC���.�݄������d� �z�8u��6��f���?Z�)����id{bզ6�.<x���d��3�d����#&��F����2��y ����Z�]5��-��҄�(
޺Y��w�z���sc�Uu��A2��j�[�a3L��*�@Nt�xԗ��f��d_y�]f~�nԹ�wt�gc�W����N�*'A����#�$-؎sG�Wj9�@+m�/�YU���,!#bB��ugjjkT���$��as2�_��YX��{��o$�WM�TL��K�bMn���*������
CY����]?\�Ѷ$���w��#K3�zR�*e�*�,�������OL�! D_m8��	'��$q��ᯁIw4�\|3Wd��o;i^��l�*��D���K����5���&sq�R�Zn��b����CМ.߸geVQ-W��1�騪�z72��V�G��ܠ%�k�{*�lY8h!@*��A�x8ŭ�xi�i��������?�x	4�((�;�j�>)�H8{h��W	�����&��W�ɽ�dG]$��>��a{f)s��q�Ӂ���,,M\��;j[��ď ��	F;�����p�'ؐ9U��a����=���|��_�bT��"F���0lwߕ0hM�Z�!���Ơc�f��[m��P���an��
��7�Y�4a��(,`U@}bΖ�h@�I�	P-��N���H	�U�}���x��Ai3;�H��u�0`pG0��4&_Y�}YƲұ�2貼�>�>�D���U�Hm}�-|gEJ\ւO�f���� y�����V�3���4<��*D�Y�F��僙� b�9�S$М;b��*�.7B�sݣۃJ6i�n��WT��_}'�ӗÂj����l��>���+�|�MF�l�7}/�C4������CcK�҃���Zb��'���e CkG�۩��p�t��Z���&/U5�u�b�"O�_o�n2,��q��r�6݁ݢ�@?o���=���~u�^@.'\���b�TeR����"5=�S���D�4��M��R�'��������5)�kk�QK�7����B[�-և>h��ԏ����]�߼�%5���H����#�$�c�<�����wK�`��G�8���3Xy5����Q���j���\Rsڤ:�V=��*��-����}��x��p�!�"R�B׫��U�p�-Z,��x|�c8&�����uԚ�c�U[[�\/S�zm�O��/��hg������L����7�Ͼ/��:��L<6�z���v1��.8j��`hF�50�ET�|Q��h{� u!M�&��g�v�g�{ς�n��m��AsV�!�ZZ�W�z�,���V�M�K�n�,J7�z�H�n�3�r���T|T�mL���y�*��0�&g�G�P
�ʟ��^u���D40P��U0N��@	c��S�B�� �0,���H�/�WG��tJV'}:��ә��F��4IQ�7�=
���GY�=�4���A9�w�A�_J�����9d��z����3�u����f��|:QFι��>Z����"�e�V�Qj_ �����NU�#U@Ͻ�]��<��wY]�gx<�Lf?�E��cT�������g>�װf���g��Z��{�t.CZ��(-�2��?jq����Za�R�ji����-�:�Z���DL)C�~O�x�ӗ��f��YU��^�@6x� ��"��2NV	����{��[�=���E�'��%�:�gDn���=�]y[ޛJ��<V��I]s�^}��rg=Ki��Q�e���3D;;;6��wLv"��C���Rd��ҤI�Z/��b����K_'T��=?��-\�U�
��P+E�<���)�Z�k��ooZ��Dh�� -宙�x�áX���sP5�4C��d��;t����v�-����/��J48��$L��G;%U���m.D�@��JC|&[֍��}N�4� ��2)���х8��M"V����G�D���n���M(�"`�(���� [R?���)}�"��2S+	S�]a۽�bY��+"�O��f`�
.�In{x)F�����BG���۲�M{$H���٘��>�qZ�&�`�eh���BSp��V"��U��r1�/ymz��؄{�^&Oɑ���̊4c��/2��jbb,�`ȉ�J�·����ɪ�b���|T	վ�k��0척�r2\Ȟ	��Ɖʄ�mԐ�1޸���=�˿�i׃)�-BU@+�a �oy*���^j���D1V)�(l�9�B���H��GƲ���-7���ֹb��0'E��i��qp|:�}�Z�IpsT�|*g�s����k�QI0¡��χ��uJ��5+.B�kNs ��2�Z��&
r�c��£!1���×!��A��A0�\s��~��-X&X��Q��(l�⣕�����u�G��c�'H�в2A<wD`Dg��(�8H��WM�V꧊8��X��e��v}�7���;���g�⡺�r�^&�j^�D9���7"fR�}�]�a����R�r
|�z��g��Rjk뱡jj+Kd"I� ���5��;	څ�¤� g`��@_�����.�����V8�i�ϝt�;g�a� F��� ሸE2�z���7��W7dN©9z�ݬ����=��C���Q�@�k!P�br�=#������D.�I�֑VF{�����ݶQM��{=��D/[T6q�@��0��	���H�4䳝sH+�	���$�	:�ձ|�|�:W���f5z�)P�1���1�w�����}��ӭ�6Jkո2,�[�b���#ؘ`.��7?�}P���G�F��d�T����8..���S\	�y�"���U��mY5��yPp��:dd�~�qfj����1�ٳG���M�4��nm}��;.���	��٠�N�0���MO!�B�`"�k��)XF`Cc�TX�Q��-����'�&D�z#"ȡ*��U	�L{�/���d�`��&��= �W�.�ӽ�ϖ*���T���Ķ$©B,1<�#9^�H�`�pJ-�_�,(h�k�;�qw�.�½��<�ր	S��6��B���[{ad�!Z�d�	�1XO�79���1�p��-
��a꿢#�T}h�G�a�mv�@���j�{: �d+¶��B�����'=)"��MuR��]������F�37w.�s�4n�1J���U">	�$ Z7Sw�#c��>0�g�tE���N������&~�D���cҞ,��[�/����_����z������Rs3v�6R�#ZE�M��V���%���M�v)�׹a�t��53sr�R&jG>l��_HoN R��|����Ťܘ�b.:��}� m�4�`P���������Y�K��S�����nZ�{�|.ေE���X�p�C�w=$�6H�qLH����5��dk&Fp@�2���v�}5Zp�	��)����!%y����u�����ĭf������LB�|7/�K���pp>&eIG(����-tWB\TA����,�Wf`3��ܬ�˜/�?��b׍��,��(��$k����(# ı���z��/�1���c����\�r@tVN�utR���|2=���'sꚣxuR��I�Iv��.X{�p£n�;���|�����܁�v�0�{>�$�Ʉ����=r*k�k�C��1���u�t�y �,cd�&ysh��������p8� v��U����[̂ Hp hȵ\1�L�ES 3��
7L��侵�����e�?^���{����������� ���������G���U�M��x+�S`>��Y����23��2��qUD칦��'��FZ�k!�6��^:���j�ũ0m��$+H4J��GʎH��!sd�H���ⳗ:��t*��_��oh�=`3��#P����� ��yJZ�k#�0W+8�8���0`��
t�U+lρ�5a����tK�L��w���7�@�s�:n�F�<]_&�o4��w%�W��T
���7H����qQ��Bb����`�~p$O��	d% �a࿓q)�){�UD�����p�h��q 86:�XDfe� �X^�Pٸ��~�G�S�f�f3d�Y������Y5���<�1�!�*~�}��L��c���O��%w�^�G�Lܰ1�&>!ZWv�@gteE��w +���L�	��"k�?s$5Q�z:	G�?�	��r�I��t��:FH���Ԅ�L7=&|��s4N�,-�C���dZ�#��<�<h(A���k�̔��K+���B��0��o�~!v�j�]4{Zy��F����L�,,&e��^�xw����u�q�0�[ih��4��&�L���s��,�� ��
�S� �շ�bT��e��(r���}�����@���\���"�'��?�Չ�؇��j���B!>��}}�?�_o��L���L�@�4���W��X��e;�]$5u-*W��*
��U��h>��Q��Zveή޵�S/�����Ow��J���������B��z���"� h��sH�si#(k�۩�Q�-u�P�4&�Y86Ȍ1C߇�ʶ�W�@�PvG�I�j�4�:LDTk��ä�`����k����}Փ�I�y_���n#���܍HaB���6�YhOw`>w������R�>�G�۶���4l���Eou���@��FR����]�BP������
�Ƞ�+���I���5�(�S,1�e��և,�z�T٣���|j���E�=�ￅoè��Qr��b=P��(���M3�sn	xP�E�4�˕��/3+����Y6�[�l��_.��&Gʥ��8sAH�m��@�7���E� �{X01�E��G~���V��u9����"9@L�)/_0���q�fh�M����I>I!�q��>8�{�VS3
���	�^?�*�>�2�j��*���y+ޓ5��2 ��I ���u���~�;1�T-e'9���,����BJh��E�,t��3S��Hsbg8���AL�ߢײ)������/m���LVrՑX.��E{w[��p���/�h"E��Ձ9�i�2�9�Y����&��.j ��{<��XL�J��R���"��;�1�EA6^Eo/���E�w�n��h+��:[$�vԬ1�'	^ �d�#�Q��u�)���ˤ��>�"�6w���7��ȝ������ӈZ��2�VX�Ǩ��{pE�՚g���'Q��*�J|hHGjΊR��D�{��(�D�
�����9�QʪN����U��ǟ����X��l�A���_[$�6��o�j5�x�;��bmK���9r���o�3�G�%��5R{\t3n?����������U��(XZ��x�����p�������c� T��r�^��&BU�b����!Y1��1���~����,����Z6�v-`�I�%Qe\+�57�����C��0�u�HڋC�?W��C]s���G��}g��� ��/D][�/���¿�$k4�`��)����0[�}=�ֶ+ϥ
n� 9l�����B�Ϻ��S�ˑ�5EuC�������AK�O�v���T~�=���h]�획ݑ�E1p^MY�֊WG}�v î��	��(}կ0��0�v4ڵO�dVB}ِ5D��T���M|�$�me��*�%8�f{�� ��������@	(,�I�K��E����|Ň_�S���߯r��0N)�|/�>��}��dR7���⒛��yli�f�'d@�<���'n�'Ոz{�f}�>B1��S"�XPu���t��곚?܉H�����1����z��&�f�G`�\���
�9⾦e��˟���]$��G�q���/m��`y
_O�*/�����?opNC�����TY�2��}x����J�8d^�8�bxS/$�6�pF�,�|j���%�OR1a����T��e�˪�� j���[�����IK���!v�F
�z{U0`�rȮ��A�MWv�+Elg��=��NAT�A�����S�Z���	t�ET� �l�u���G�1���҉�:��t~�M�7T�5j4e[�e�=E*������:@l�c.U��$}�&�gb����U'�m�����
��7��I,GfS�BgSN�JI�rȓĥX�HӺRD&�Lc8h?���t<Jc�+���pږg|"D�&8�/CE)R5�<x� ���c�Oo��򏸅�U�x�Fz�ĊC3u��^�ߚU��8m���n�u�~ff�os�9)�����*������ǽEL����J�y{�"��8���
sJ�j�{�����y�M�ȷi��/��4��fi��]���g:#���Oh,J㰑��ݹU�1��m�᪞��'��}4@���U��tF�c���;�mٞ����ٞFQjE�,��BѴYe<[��H꼉��U�E�$6��;��m�r��/��=\��&�ZA���%G�E��̧�z�����^}>Q�������$�_0��Mڄ����5\�����Zb���:��^M��*a�٤�B�^6�'q�x�:�On3M��S8����������u��j����8�D��+����-? �&�tSUq9s����1�!�����iEPH-�4���iY'*����.�����%����X�z��f�D͂�^$S��@��ysBQ��t���1Z�r[aͫ����H���H78fm��"l���i�"��#�Q����D��%0Z�v�ʞxщ��.Ǹ�d1��,���i�Ǹ0�hNQ�T>�\���8�&kB�0��^ܡrH�Ԥ�{���ه-@}�<2f�*H�l/�ng^
0�Qd���Q"r��ċ�L����JhuX�@�RA<z��F��!�|J|���%��
�Q;lN��%�5��0�z+�q��x����3��ƴ&8��d�Vm&v�����'�F��g�Ѓ�{��o�b~q�p��^�tu� �_�ߧ�WXn����!6��2���8���R�<�QK��]]B}A�b�6�HG��*�<��O{���{H�W���שR$'���Gx�ʝ��U��3v~�Q��r�]Zcp�<��1�����Ń�B���T$�:i8��@����6��l%Z���M����ԃ���&���Yⅲ$�3
�W-k��.׌I�:��|�rZ���w|�U��/LQ����� r^x^��7��<�z�Y�>�
�ro��4�T����F83�.�r�{"��0W�0��${����b���ۭ�3fgc�k��L:I~�����U䰞Ĳ�h>_����P"���.L�w�UF�y,%v�@<#�>\��w-_��W�PE��7#g��㺕��eF�.�<kT�:��E��p<��x6a��Ҩ^O���\��G��9���K('$�F��<���X �g�:VK����ԋ{tL�x��V?V�_,���%��-)�mP-��[GGԁ ��d<n;C����L�_&�=��e��0i��Rp�f8U��{I��x5����9��G�,�ןD$+2oJ�+ξ��?�,��t���B�LL�#������(L-}�CEJ>��9���<�$Xo«ٔޚ��ܶ�v|���{u8h,����ӰO-�OiBp��!j�����'�D�@>i������nL�Fw);�<�_��ce�S��o����&]�]>��ו�w��G���H:���ݔ�Umu*�о���<;�M4����B8�f��T��Z�����T/�BB��\E�nJ�G�MU�9I����Z���"�ذ(�G�A��u�G�A���I�iRH_�����J{�&��[�����E�� 5�y���L͸tL'�9ٓ������#�����M%u_}�f@��nUW6�y���*�\s����54�G���[� �� 'hq2�>�7I��NV�.�z�������Zw1qL2��T�q�\]�Nu�%R$:b]��Tm#�ik�8��S>�~(�$�� ��(�:�������{^\��qK6���FY+�i��5��A�؛D����H`}5QH[�p��O�Q�w�z��*�{46k&�>T`����i�eI�%�z�jH�|�)�ְ�46�������LI��Q�eIA!W-���U���W0��]�C<�e��Lf4jď��93����1�\��(�p� �%�Ӫ2?�Ie�����t$���~���;8���r�f����GU���É��&NxQ\�\K�tK��8NOO��|ń�I�^H��lS���qbБ����û�n'ˇ�	�`�L�e�zuqD)��w4v�0D�GBAG���]R��	ѯX=��ؕ�����ˡօ�}Y4عQ�ж�P��2qv�i��m�:�8��7C�p���g����0�Ltt"�J����x��ُ������R�8��g~dȒ������+FZhM@j=k��q��t͉~9�W���"t"_��m�KV�r�QA�#�'�e����X�qH<UB\��F?nә�aB���Z�'��,+P>�h��nZ�څO�����5t���4c��?/A�L^nЖ���mp��V���,�u%�@��
��o��Q>Z�JbQm�df寽Ư����i�/�#��O��Є�^r6���K�UF�E�@��PB�Ag�����h(w���*R���߷l5�_�Os����½��#�b,vz�6�3\H�eL�X�mMY�Q:�"V�J@]!$"�q�>$�r��6��u�@��2����Jm��{�0��o*�@RHA��u*O��k��>���*`T�s�"�9r�Qdg�����wn�(�@+�EaR�V�����ἑP7�hWA.��)�s�ha�+�;��`")�]>��3e� h|���/�*�"y���J���?�
%_3��
�����׻����A\�����p<�S4ؖMf*�;&��nb+o�c�zF��cF����O	)�6"%Z�8�Me�&^����C��0F��%$�y5#�;�bdc����c秮L�W΢�dT��ARv���#�}�:}�+p���೽ׇ��'IX�����a8�7Bm��P�mW�E|�t
V��o��ݺoI�D���O�����_�OU'�js��j������O�)��d��krH$S��C̖������7D�f"O��~j��������Tp�+�GH�C2]H���_c�����	�k^ȹ�f�ܛ}���䍰��rƕ��W�[�ƌ&$(p(p=js� �jM��1�Js3
q�鲃�o���|��jNbg��Z�	b+�N�e�Ձ1�\ī,�s����UL�f��io�Gv"ϓ�z��1jJu�nժ�-��]�-h���@�H�UR���α(c�����%������T�ǲ{�M2!�Pa��T�Ou��N����fr��28qu gzBg_��+�`[};�ѻ��_��v���4����|�^53�o��ģ�N,�c�6f��B��Y��?q�X�HU����"�\6@;�ٝ�9�{=I��)	n��ɨ�� �.!���v��|l)�n��wgڢu+����ƻ��z�!TA,U�4O�*\�2!(��������[�Y���\[w]�Rc<z�� ��u�?�/�V�phLeKEU��]�/Vv�/���O�e���
)Ű�.�>����4Fg�e�V�Q~WCd@g�W���㕾:f}��q��
����t�5UX��_��O�ݙ��Œp2�%4�4��TQC�^����ʕ��k�җ#ϱ�m~(��O��x�{a�U��,`�~�m
* :t~dt(فʤ��:�~jD4��n:�Jv��7 �����Y �ܜ�r����Z!�y��ٷzˡ?��m�Z�X v�`�^̉��ȯ�mf0��=*a+F)���V��o3^,�;X��W�	Eӗ�{;������Y�O��wA��h[%WN^پ�$#��*�y�u>��AA����,(p��'�@�va�	u�އ�!>�cuCR<��E�-J-
d_�љ���
<p��&e؁�&�����\ՓFa^}n�O��*k��Z�A���d�����J�"�N���䝰X�2�cԵ��br�&�����>A���@e󐄙�>+�ʁě8
��z1�	�uȽ]k��f�n���?�P���Q[���'ß��Ŝ8ڃ.q��|N[�Z]�T�����SH�!���٭b-BG�����)�U'J"Eꁡ��Ѕ�����6�\܉I���5}<�(`r�K��\t_"�5���v��!4��.�#���.���4��F�d2�v2�w�O�#�aqܫtA�0*�;�;�	���h*��ӳ��8�9F��q���?�h��ꘜeeY��X>��7�*,'��̠���x���?����������{!��$)�H��8鎛�'tX��l�n^ ���~�q�G���=�����F���鄿Qs��v	����W�I���F�`ƪ!#5jM��:A����)�[x1 ��.�������������g#A���@+���Lk.����b�tK��U�oV�����"�h�)��*��NV���SA���>�=ci�W��\�K%�0��@Kpn{�ֱ%��t%�}8�Q'�h:I�i.����n:�0V�E>������M����g1Qvn�
/*c���ɐ��,{��ei���ڲ��(��(CP�k�Cd�:��0_*{�����B�w�fz�Ϝ.}/0�5E�� '�9X�X�5y�6�;�0�w����7��_}a%>I�6L������d��|����u�(����Zu�}�	_w%�ؘ$�L���&N8Y��;t���ݛ�N�$3�/E _#�W�[3F�]6�Ƈ/�����+ؓ@Έ1t���>B|7h�ۥxM�+������٣��2��d����3Y�it�#�ŗo��K>c�;2��������j��&gK��03�+�����bR�%�]�Zz�rS;���&4� Af�+��uЪ�P
���S���۞& aK����������e蟁���Ka@�]}cRzp��`2�kvu�\p$��о�%�e/<�5��lFS��Ux�`����%�Je�k��b*��󿒖��J�Z��Lr�.$"b17��5z���9�����2Z
d
r� m:������&��3�qm�{�F�����|eaT:�YX4�"J����n�]�CM��9#v��.��q*%H�5Q6�Tn�ۓUz6)��-#�R@o�c�82�5���Au��6������!RD��H��5E������#��G�+�c
h����/�6qW���7+@�1m�R���Fk�`��<���H��9�w>�Y7�1S͝G;����s��n��@���� ��N�yz10��4��|�֥"��?\�İ���=4���K�M6؁�/�Q�R�m-��v�5�m�,���
��2���L7L�˶�:}�MN;���IZ�V��eM,�!t�T�I(7�|�oJCl�Fl�%g}���!��_꼴�
M�StJ�D�U��w�2�@��ǐ�	T1W3���{�������������"ՔS��
��vho�W�vk��%�Ϣ�!;���!r��.��A�>�Ԧ�s�׸s�jP�I3�$ 4Tt���ˢtr�W���U��SEKh�@"=��O����BTE�OyycV������9h��W�~'4�;�8��T���~��䱰/G�v��ۖ��$W	�o�{9�j�X��w��{�ZǦ#}q���5��a��$d��7�^�Z��g�&b�zv�/|�o������M%��\T!y�p@�nL-E�k����h־�EG�q�,
p��C�Z*":[Y��,qJ��:,ix(�3<D�p�5kik�h��'k�yo!�V�	������33��
њ�C$�x3 �-�ݛ�ZQ���5v���ǯW���}���D|���s	���L����{�+���	Q(��>��&��p��E�).X�����v�A��tHQ\����CK����"_���VS�S��z��c���j��ȶL�M�?vj�T��Y�t��R*v8��|)_}]�9r�ð���ѹ�"�᪬�V�n�\+��ȑvBH��;��5״�t�Cq>��H~����(�ֲy�i�ǫѸ��QX�J�W��c� ���|�� g'{y:>�O� mc��ƃ�)ρ�J�D����-�}��!����4t����$�w�~fg�0��l%�q�h_)\Yuନ\gkھn�����N
���9�� S�K_ʝy6w���L���b�>������2�h[_5����@+��tD��HW���v�0rz0L�ܴ�4b��f�Xi��}ŝB��ww��d������6h�,;?��4�?�ZB��u�'n��r/.5p̙'wb��Y���A�u�z�T6�u-�[�@|!�z�lL��<��P��3�c�}F�&_��>뭐	e�ޢ�$z�S�Ru��拍�v�Av)qA�y|i�ꂢ��qT��a}|��E�?oп�+Io����B��I�z!j�YY�[�&(dI�Xp����O��n7�t��Ϸ�$�?�ai�� ޒc����mŏ���Cz����o�h��b�C,�^��_��x���m-N���SY���V�>��(�߿���1���M"%bZ�+����y="-B�����*U�fbI\�V�X~5�dav�0(�k�5l��C�6ĉޒ����柘��flTJ���^58�bj)�����ef�4�r�C�՟<������y��<R��`�)r�����	�P�e`�Jp�%���i��>���mT�]�D �O�x�~�o��R	5c$	3��fd1���Ͷ�s��T&?-nX0���d���x�U�ϫ�Xu6q \��~UW1&����ߒ��ܲ����ۅ�����Or2_�ۥ�%3�7�a+X�Lz��9cv��6'�CSdj�����=��߾X����~/�dpw�m�aK�o���+�����YQ��d��f"耉��CO�k����ǐ������S�h��@c��է�B�x4!��	�2�`���[��Y����3Q&BT��"���9R�E �{��m�d{�������^A���M��9�`~�wA����/醾���,DS�B)���tYd�G�Iܥ��ꛌy7��Dcs��}{��_�G�gI%�����uQJ�����5b�n��)eǖ�����ڞTR�b0LLDЏC�Ggc&C��ar�R�o��H��.Z.P�`Z��C"�g:�~������7���3�N��R	|��x�8X%�1&���O�6Z�[�0��5r,��pe	���=��bs���;F%d�e�I�(���"d����G}��J+&���7u.�>Ȕ
��P+��]��D���b�C�ɰ�	��ӫ@��"RP�j}�(i�G�?�Y-�%��N����d��?�!��d	��B�����l�����4)��MC;M��T^�ٳ_al9��u}��%C��i4�����uv����r��o�,�7!U�6�!�Yp��OU�=��~<�i:2�T�p(��(�;�m�(��=pc�Z�F���I:�J�n��L�8�!A�Y����"jx�.=C���>���Ky��*���W�5���l���{�!Ǆ��7sO���k�M���Y�va-ޠc����酝;�yٿö��í��ɖsU�> �!{�[qo
�U�!���b(�.�еhc�Zxe��+he\F�U��X׹#�eO[�3 RJhq��2�O������V=�L�,�1FrܦDD3�� �t>��y��X!�a=�c6�i�"6%��2���j���U��(&|=M&���4���/쬟��  :ň�r��}�?���� ,�nDd�?�!ќݭ틥��a�Xn�`���2�X})�̆~��̘rbĥاK.���:���,���N7�\`���l�RP���b\���ިPC�bd���D�����|�6��b��&~���	�H׹�a	}	d�\2�����EY�x�.�W������EFmW�[����ɷq��_�7z��3�כl-a���1�Wl,yۆ�iJ�t"t��%j2v�MHL�� ����5Ue�-�sr'.%��^���*�8(�J �w�/:�����Fo�x��討�J��H��3P��7D[�4�M���LZ�M8{��~�]�J �G�,%�r� ��h�C�w�z��8a�y���vQ@|u,6��A=:�TIV�K���↮����n^���5��"�Kq�����'��`��x P�4�6�rS< ŉg�(�A��`��zGu�� ���NX���0D���x#\x��r�!��bЉ�Ь�T_+964r��Ѹ�����tvia�7�'4�U��8",+4NǊe��x?펬+�`�6� �]�r1}���Z��Ă6,fR�GĆZ���sr��E���5	B�<�G�9f��K��<<Ew F��r2�.�|��U��+
�
��ߝ��5�b�=��9�
5\��,�+�hV��%:G$�z(��BV��)a���v\̶pVFg��	M�y�<��ǾC�����Ր4��� ���+�ϕ{�i-k�+N�،љ�Z�c��Q��Q+v5k[7iz$MC���I���?�]T��'��.յf�̚��rf�+��3�m��� ���$�ܾA.S�M�2s�*���h�C�jQ��Q�H�Ix�Y�6��Li�ڻ�φ�EU���t�l��Λ�D�y̓��AX�ZZ�6�"-�{+�4g7��u�4hxU��s�P��n�٥M�f���f�#K�V�kL���aQ��~\����|�����٭zb��I�?�ک�sv��p�6K��vc^FY	!�"b5�Y~�l��q���y<��na���g\��ͼ���v��Ɓ�0�9�W8?�@�B��}$����/���*�\��/����W]����7�3�.u��
��J�#n��4������(_���mL��W��c�^�ty�B��k�����2��r{��.����F��$�R�X~y;��O�����e��~2�/fbb�n���3���P����ۈ���Ya�g�T�8�=��-:@-K�Tp��!TZ�����"�:�����(�͎�m2<��ëa��oĞ�(��5���f�.�;LD��	�h:�\`*�&w��ɛ��C���l��C#��D���h�J����])]J��E?��g��_y��H=���5SRYG��3�M��v�M���
�R�٥�L�
.��B�V�~��l<�"���F�kNmngӌ�ysLO�i�¶N�J�r[��q�豨��@Xk#%�X���r���4�ڕ�0��p
~���	�����@]FiK��<L�V�_����X���_�����,��oF�r! Oes�_�Ҁ�P�2"�_ܑ�U�ܫm�x�lN�l����0J���i*�&"�ļ�����f�ע��#��
0=e&4
����%��p�+��)t��X�_��r�[�kH���_'�_Y�� .SKψS�R��l������kX���t]`�%X:�訣�5�HQ�"��$�yn/4K�<��F��9~�ई�uE7�~�#�uh$0i&6�μ�b�3Z]'��S55��/�@�
�	y'�e�O�xt9�s'��y
�# ��u�	�7w���"���ط��װ b�P�/P�[���"&֯3��	�����T����ax�Y����m�D���ې!�?��d���:Q4��K���v�{"�߳>:رϢF����g
G���~�;�eC<:,;��b����&�d9���D(Yu���H�MLL[���P�/X}E��_��d�Ў��]3H]?�oUX4��*/m:���Cw��ۧ1$Z(��M5�f��h(l�O�����ʐ7(���s��-���6�O��ʁkkF�2�:D�V���aB�j��~m���W�T� ��$�j�<�d��R�[��u���B�P=�Ue�;N�:����嵼���G��߃dm�M��������s�!��tD>��v��GW�؉O�/.�J��n�ׯA��)��:����Lp ��D��H�����s��i�<�LV'Q�'�?�'#�O���w��A�2�����������m{��r��ډ��#Õ�W���g�0O4��l�"	�ѕ#<^�"��Fw��o��b���~ �g��F�ǇJ�c�}���;+��|D�O�-��$���0���U�Fa�i��j�DI�c?Tz4���LJ}���4���T:�����`u;G�!v�ũ�1�\v	��Jdd:�A4��� [�x)��/�9tjB��Bo�q�� I+ā���A=��E�>����E��~�;�Zz������u���a@YѮ;�M���\�B�jn��K��^��v$��M|�K��ӛ��q��]��h�y��e[
?a�U��dW�<�C��P7-a��V+�Y*|
�@��4p��8���;�wR^�*И�&�H�6y��5�J|Xɤ��/ӚEE�[ȇ�=�8<������dz��>8Bc.hf]��ʜ�j��,Q��������1ߟ*���U�G��:I���Q*ք9َf͝z���0$*�?���'/҂�O]m�bd��XMS;#�/_��G5�F2�e�<¨���IKT3s��<��nb�=+[���o�8�d`���Uy�|{WY>���)a��`ykN�+X| !��̣�G�WBM���4��]QVo�i���)����5Q�N�A��4�xk	G��Vs�`���mS6�sm�#�*����1d ��G^�Ѹz�$�2o�m���1�Q�5�ؘ����`�I��aE�~�D/�U%��?{^��h�`�]>NӇ�e�I%<#�W�mpu�9�+�9$���eX���ke�}��s����-�aqlYS����6���?P<]�1D��f�6�N����D����a��z���/=�Ȭ�PYV8��q7@�oN�Ƒ�XץU���_���X#�b�̺���iR�M�<g*���?�lM�����$y%`~��B�c���B� ��W�:x��P�[�QT��d��b��#0{����;:wO�jÅvl��Un�wk��+�xB���v�~�?�P�F�/02��k��̾2۵-Cs	��|��ӗ������6�Xp�S`M��_��L`q�1*�M�Q��@�b�O2(:W�������������Թ��6�Tb:��I�U_����]��Вa�0{�TQ���%l\�����P����PjL�HU�������'R�"���շ���Wac��BdXz��Q�� o�Q/;[����Z�����$(�=���ێ~�|A��CZ��.q�r����[����ݨ��A�����Ѭ%�{-߫�-eJ)�ÃT���G���a�@�#W�'���o>޴�
���:��, �$|�s/Sb���`��-�6sC�I��i
m�t��6Wu���U��̍L�e�����㿿ړ6���R�M��X��*�mj������\s�y�h�����-4܃���D�1J˄���a�M!�0r�oJQ��Y4�1�gX�x��J\�R�EY���� e��v�Kz�Y��>�ZT���i-y�w��II���s����^��'�(���'��o)���{��$'��v��/���_1 �w͒t��ƕ(1���M���ɑ�V��{��v��s��tRP��[�	mc����ѹs�\G���R�p2��!7���͡����??S�A��h�}697�]�s�s�CcO�3���l�UB�!E��姠*۪9jr������ُU�b�v���Y��V-QY��#��mfG*F�j}��n̫V&=�����`BW����
#�����鶫5c|DF'�0�괲������!6)jw$�B��AZa�̂�K���9e�@�mw������(�7'���<#vn!�L���OӸ}�w�w�P̞{����� ��#q�5��r���o�^Y�Ip�J.�?��GM�el(�qG��_E�;�������.M[����m�S�qAۋ.�s��{�:�q}:hǪ�٪���dE������ �o$��(5σ���m?Q��W�g�.��S�����>L褦�+.���;�#z%t�5R��C�[rb�f�����<�(��]�
��C�x���Z��&4\����M�13F���	��#��`I�iQ�����Y�qXDO`�R<X�N�dW��o��2 ���&�$�04N���랑��\t,^/&��SXk��:�Mo�c�3��5S߹Ȝ��s��U�����h�Ep1�]ov[�̂��qYD�:g��*�a�S�����~ߋ�gJ�_�:%
İ|"�Z��T��Ap!��>U�5@�r�����1C�hse*^e�>���{��fixT���滬�#yG��"n@�vU����d��5�.MG��n�*r��"���E�Bs!Έ�ne�3���a���塲[�1�-3gt����ءO���.�<������Q���_QQ�^��kVD+���tNF�zжI�NA~`?"f�����9M�X��ʅaUg>;�2$� ���}nǃYyt�3J��`2���SN�*�c�_{��|ߗ�~������d��j��_NA&mSO7�r���g��u&�y����
F�&8ʈ�2��w�h�O3é�r>��DIT~�əB��Ȩ�2L���뫀������ml/SvEf"��٧�"���:`>�(�	w8Y�A�TqZ�
��7�*&���ߞ�PƱ-��:��賛U���R��+@QF�mV�>��G�Y/���P��/�}�����4��2udb�䧴���AFP5�J�׊s��Μ��'�;-�F�V���b�nV�&~*�M į�O��K[�����Cr�fa'r�+7%����)���X_�&{AI$W���?F'����Z�!׉� |0)v8��,�Шؓ�g�u�n8���2{5XZ�]�����4 �⤱y�����ϴU���:b�\Ia�dƪ�Ûby�4g���T�F��ذP+��lA���H��plWB)��4�;���̲�+\7x�}D2�w�� �ˀ�w� K�����˻��&��_���֭%f�9S	'���mA�L��Zc�P���ZQ�m�?Q�Vg�J��̀�b ��v�뉾M�x�E2�5FD_��ʪm,49 !V��BfZ�J���G�X_o�wV�nX�Cg�۽ F�/ȡ©�_+�+3�тmש�R����\�����1��M.P]�o���[��q�s�3]��݆b�z���9- �P؝�,�����<�da�1w��qgd���ӅL��JyE�Q7]�{�«�v �/R8ݛw��vk��6�I����q̰(�׹��VD���1vm��FC�Iz6V�Q6邾+�ʰ?�m>��BDFܭB����p�g�6�H�>n��W���t�� .�p�2�KrO�����2��.k�y�р��:���@�����E�%0��6�~�0����3������f��o,���Y��u��--~aa.����U����;Z�c9�Y�-/����oA�Z{5�m�.,P~Y0}l�D��uN��m�q+�����£�ڭ�'��.�k���򫍔�8o�{�E&�L�[
�iZ�'�����>SN�@�Dx-����U��#Z	t��^�� W� �}�S��][H;$c��r�}b^�&��h����sfx�6Kp����+.��׾D�~w�z˔%�~q�c�1е����#!!)�ގ�<˚L�YV�����>H`���m\7��m��"��|��;4��b��I�����Qݫ�rn��V���PoN���{���ULq0V�\G�=�*��L�*h����Ӛ��Ry"��g�	cUO�/�A������3b�U��qG=�c�U����mL{� ��^0C��r��^��v�����͏])I
j+T�ϫj�o������Q����H�Gڢ�
�_	�,�0�'\��������<�E���Z{
��ߒ�x�Z{h�F1Š��:*�.����=Q��\{fC��AIGVK��"Ֆ�qe��EӴ��,����o��)���|FBI����c�b��;�w�j�1���siH>���ۆ���Ȝ��;+
�Vn��2��e���0��Xk�'�r��m�u0�4�����^��X�)�yW�k]V��z �U���	�Fg�&��p���ev��ϮL��~nC���K�����;�҇��.bĖ�2�ڷU�-%%q���?�{�&�F� �up;��	p�(4 ����j{Y����Y���xu�:*z��7X�:B�f�r|�UЦ�q�C{�̼�
]��TA�;�LF[G)G�v J�=����~z==��G$c׃?��˼l�U�e������]��2n�E����q�d�K�3�U'7�D�r�(
�������C�J��ZI�踈��aڟ��,g��)��
��0.��%����nWAvl�P1�TI+���#�	����f���J?R2��@pV��ӕ�}t�Ƕ�0} Lal< 2�y��nmЌ��T5ks�W8� ����4{��44*��:����7{�;��	�	\f�VB.�X�����bl�Hhc�n��l�O�)G>·�#2�۶R�?�M����:Ғ|ۯߨ��@�I^"{���]lv��6����u��V�4M��9� Jz�?�a��_��Cz����f�͹@�aWn���*��حr��ւCAWk�������Kt�_w=z?z�T7�,�ĜKŵ��K�sb1t$��7	�ﻥBPs��f;�"���R'���J�M����W�pYߪ�<��+K$�����~9Dp�����Y���F���ýyS�Դs����W%	++P�o��r�n=��DB�n�����7ZK�;0�^l�w��Z��H6�E��(�_�3�� Y�Bx-.���nm"x��aŪƝLw���>��MB`Ѡ蝘�_�����01m�j�$�~QǙ�$׈视)Z3]���&���,�����"v�1�����w�!�=�Pv�<��fF�ɒ^�@��#���E�ɟ�Z����2\����w�Q!-��������������G���/�t�,���\"���G���>���j�el�}4"~	ޭ kw�_����f�#����N���a@�����F9?��2�i��S��G6���u#{��dxF; ��bɩV���ѩ����#}��c�p�[( �4Hj�k8^B�1�t�� zt�w�p��L-��_��bI[��E^�~'�$Y�_�*=����,��Σz�pvʻ92K��H�}�@��SJ���-�&�:'�j(�oQiTg�#����v�I�.��/I���&�VÍC H��-pY�^u�Y^Y�O�*�/�ς��*�8RstWaR�tb~�qÓ~���i�y�}�
�F)�ǿ'��b�]�l��_#1ŗJ�ԇ�##֤�Ug�8�'��d��w�\��9׃~55�VA���>E5k���~b�n�*�g����R]?P��?�1r	ޘ�c���\Ձ0�F�p���&ڶd�pѧ�����}��=!�����y]�J+27����@��E���I��\�^���Oz��Z*��0ǚ���)���[�a�B.�R�"�*�e������1��J��c�=�Q��gk��B��Ծ��xoZ?���<^ղM�پ[��	|[�h�֙�A	/3c&��ݲq� sӇjĘp�D��ݍ���C�7͵���6��KCJ(��ɣ���f�3�	�F(��^���F���:Ա;�HB.�`q~.+F��]q֗�s�rD��������]�;y[�z{ ��0���б�"����Ł����
bD]�Ԑ��������7��͓�ޞh$��z���3i3�ɿ7M4O��2�<�*+����ID��`͉����,�S��3�<��E	��x��$3�����qB��ΈbV��ϗu�#+[������KVa��#��ؾ�����_^�J�b���R8.
�O���S8ūɴn�LP;AW�A��9����o�@cP��K��+��F�N?�Ƶ�N�y���YEޚ���;s!�����+�b2�I1����k� ��(lB�i2����� ��Q�:�~�_��k�X����D�w$l�b���UQ�)����c�S~%
��Bh_^vhD�H+E��o������&��=Ⱦ�~�*���f�;�1]�}��֍у
�ɹ�>�W����I��X�.��6�]�ʫ�^���}�]9�9d5�ˊ�+���A7��~��pwhs��хD�V��F��O���z�@�g��#M������Dˈ���2{=-�;�V4h�Sy�R��>�|!�Xs}pJ��ꛌ߱6a�q:r��g�唀 RX�i)�g�W�r$;�!�,�G��0Q�Ϻ�?@�����|�+�m����B�F)��V_^H�p���-kѹwf�;����-�I�Y�12��{�3p_� ��|�,g���8l�k�Ӹ��Hi\��a56�8o�N,)�}�$&�^� ��Κ :�2;��K�Mn���'�����ԁc>����(����5r��?�sۍ��H~@��iƐ3MaQǤT������3��R���X��F�MT��'�(4A�i+�](IkI�ry�5�M�YK�Y;�*p�_0�t�T�/6�NĜ� u�OHi7�F 4̗���5���RBp�W��"2��NA���O������;����@"o�k�d��K�tgc~T�hv�š{�Bq=��J� �$�~z$��r{�۶�E��Y�L��P"�)����F�:O���0\�k_Ŧ� $F��F�pG���8j��ȶ_���%�rS���8����Ǎ��?�,>�Ĳ��7�N����N6b��1��[Y̍��n�4��������Em�o��l��@%:��	.'�>Qe^ɼ	7��%�}�O0� ���Ό�@�c�6����;-N#��� 0]k�0�\Ǜ;�X:ڃ�������XZ�x�a��-H�΂��\���)�Ǖ�L���*O_b��z{D[�0N��E���c��i�>�wн_�{\�pX�S���|#!��YQ�P�1�
����0��zF-ύL���B���5)�"ֹ�H�%���z%���|Xa�yEJz��)a`wE�ux
�U0o�i��Z�R#7v^-@�5���V�3�W�%��/U��듁Bn����*�ٍC*�sg�7]J5s�܆�
���`��8�R�W#�>^�Gp����O�5ՙ{�g��RU�p�(FSE��<��S�	��a���!~)�c���.ڶT����3�|dD���`�����7fX\_۠�����1]� PN�ῆi:^���:� m��d��p���sMO)v��L lW��Y�N���;Z٭G�s�Ӆ�'R?��I���9����pź�4�c�&�T�� �����1=�ӗx��o6U�p�!GI=�t�m>�m���߅_��>C��QVrR�+a�������Hv���"��@�[�p�RB3��vG-���J��A.�'gsK�IYZ<|�wR`�*ZQi�sʥxO�����*�zn�lGl0�0�5�&sIv)U��Ý,��<b[CjY�f�DdSZZ��+���2�����U`�{5s�={>��nj���ǅ�+0N��bF���gb��T<`֭,�BG�Ҋ���q��G�`�j�"����������3o*���<��V�n�&�u��0��yd [���]���i��`�RDW�=�?����s}���tQ.�R���c98i���AW�P3����sfS�c��FY*���/���\������LE���ѽ��2r֑�z��2�ӓ�\�F��а���a�
��L|O�[���"&d����B�*׉
�^���@�G1 �۳>`�f�:�&[�6JMZ���QX=�W��*�JI��(�����F�����q�����"=ͩ��:k<�gܲ�b�P�|%����5+�N�Z�$�$J�#����3QG�� _�I�:#�~��b�ˍ�YP{q9��Jϴb���&?ӹ�M���a�]n��K.099��0O4���%�ǦJ�0�/��;����Gu��?��X/�dha�re5�]$���.)�n#�2N�<����
��H�����*A������C�����0���Ikc�'t.��yG���`������)�X(�px�irsELFEω�"��nD���#;�t�I�3gU�HtH?�6��J{��[�|�x�Ar˧9��;Ӣ�)%�?ĳ�e5�����|�����Fw̕ȏ�>L����:+lΓ8�x@�O$ӿ��Z� F�Y»�'�h�=�F��3�	��J�C�RB���T*+�(.�:U��*l15��>Iō���I{fc[�\�k��v_����A��Wp�4e�|��[Q�W�R�����|c�3u&֚(�e����(`���鶚�����.-&BO�Df��$1g��k����|�|2���+�8��_��埒Uw��O٫��P�MI�$H:	Im�z�_��3��dJ�|���T�2��o��or���D��\���z���Gb���V�;&�O��m`,��k��=6[���gn ���ѳ�~�^���q�zQ�<-�29�6&`�z-o6!�n��9?Ɓ�)��:����f'W���K���9a�?k�(�m���� ��s
99�=�dU�q�hca�q��pE��ig�T"F�W*� Ꮅ2^�3&��W!k͑$�{j���Ũ)@m�� '�#1
v�f�q�F>����[����� ���u���(L��4Ղ����<�bV��&��TG�ǵ+Z��b���\�<GK���_t�f뜔�L��ĔjWl	I��JgGg幒������f
�c]�46@��	e��
��% ���+����зض^&حJ�'&(�5s�3FꙂ_q� �8�j7��L+�]N!w�#QL�Bާ!��|�G�	�dl�-A+[L���SM����o����1Қ �/�¾�K㡧��V���2O60pa���V%�㭡��H���4�ћ�GkX���8��|��%o�x���`��^��tw w���`��t� ���ְ�����ɧ�T��~CӋ��w
�;j#���);L�O:��R2[�G��%h�l��<�(��TOɌ�$/1��U�u����z+�-����d����'�c/��T���kJZ�܁�F#���$�NNW�/�
8댝X�16��R�M_�)��8��(�,��A����&.j�
>�x���qYJ2�ɟ�P����+h`�-;�"��A��������������T�7o�9~�r�0�����A�k J�x�TJ������;lB8}�u�{�X���R�/�
y��Bp��UF��Z8���U��p|��NN �O������D�"��#�`�t�B[�O�F�ͫ����|��#�W���1�����1�C��k:ߨ9���ۦD��ws�P�a�r��W�5�*?�L �ڂ��3H'��O�9��U}Q"�D!���&��mex�hF�*(ҳ���%�x�Q�8�;Q�8�/�BO�z�m�p�g�1C�v/IgH`�5Mp �po�s�bܟ%�yB@�o��^��]��~�U瘻�{��g���$\��
5��.W�e� �[�y@�#�[%�s{p	'�_�u��Z�f�Х<�OH^P~)e�N1d��q��M���q�L�6��Z��3=!��[��O��a������h��Rck��oN�W;O�Y��5ۣ���]�p�џ�x*᳨6n�p��ݘeMe�[G&��<���^��(�.>;��_n��|�$Iܯ8���(�	�#��n7����qgu��b��;��%	��j�4�xeA�ҽ�#��SQ�(�2�Ȇ�l��:�~�x1�@�� ����;��~	�<�����	$	� /�x���N"�7��JI��,܌.�N�9B;c`TW�DO��Vg`E�Y�9���Y=�'��Bbs�B/ڜ�fO9��Ϋ�6��3V�$���z��y�y
�e&��Vk��t�X��t�5��������3�8���>���1��rCh{��?�¡m�I��I�����j�ŗ��h�F�(Kt����#���?8U*�c��YY�r&gN�\l��\��.,�b�*|��j���4��s����9=S%!r����UG�F}p�zp���8|9|8�q6��M����D��������-�T���#��1�	��� ���V"3Td%�<��[vX�^��2iT�W:�T(�˒6�����Z�1�?�GmM��u�R�6H��bP��SWد1����?�}��~H��%{1e
!BT�!V�J����jY����⼆��g��t�L�\��i:'x�_�+ ���s:�6&����@��xf�����۶���_ِ�?j��&�+��s���� �r�W�H JD���F&�j<|ĩ���8=\T�����8��,�z�v��=�n��gH.BAJ���9��E�Hɚ ����[L����(����,�{E��5I�/��9�7�
����������TVbg�qu�B��|>m2g��,�������[��ȴo*�/�;�$
'-�ǛܕW>��mkm��g�,���%���]�[� q��Z�xt���
҅1J���(������l�J�v�����n��U����m˂�Nb�"��b�(��G��k�����Gn��Ѧ�������*_���J�̐Ŋ�f|"�=�m{�SR�o�ӅD�|����zq�\��2jR��zA�G��)��	��0�
�A�x�g�<ߵ���R���δ�\��ګ���*R2�b����)Ĥ3��T�Ŝ;#<�#�g�����DY4���E�ؘ(HJ�>�TO��<@��2O�	w)	������<"���3&H�ej���Q���1O�������i�U�C�������h�����B�\��3���;i�ϢRx���J*�ai��b���v�ND�E� ?�n��v.MoDx�I{k[�u���xĪ3ʟm�lz�����.hZ4�xbn��kz=?K��(�ӡ����i��ǖ����%�ho�4�Ȟ�b�쓁�"�T��E�Ai�cin�|	X�'PTL�1;���y:�ɚK�FO;{��"�"�}m��@2�����a���\u#t��o#��k�����NH�����HW��$�&lw(%�As�(/�)��3�:gU��l�q�Y$5�%^��{��ޜQ�N���sT�5Ift���wB�n�H��a(���M���:��9���(�Y8�)1A�="=r�,���?�KU3��@N��8\����ʹԴ�l4��v�H7�_\,��#��m>�L�����	 n���к��BI8���Z�3��|[L^n0�>h���V^OV-5�y��o:��$�����Ⱥ�9����LuZ7����M���.}����JI�T�l�_��Њ��_>�4�
�߄&#��5�OUZ��@7�8�X�U�k��Ke��H�C��l'e
�z�<<S���������_ٟZ0R���Iǭ�#��	�L[�u��p����H��1(=��$���� �끙�6~�0��ͦ80�@D�wkf��>�R�fS�~����4�t����{���4_��'�9F~iu����K���XP�f6�����^6�F0�+:�sw���������Z��"�DRd����Xpw��Yv�J.�����NL�H|�(��	�+�l���>�k�0o�z�1h�o�������*��6��$�]O8
&���8O!�X�랆��s&�*��D���R���������."����Q;V���\Ks;��w�]&|��@�aQs��8���v��RH�h�G���')k�k���PJ�Q��69Z����dL+�0�] ��bRf>�Fp��� �:g?��U�|��y[X��R�"nh|Q�o�$��76$1:�Ɓӭ�Y��{<�4	�"X��D{�ϳ�%��j�����Q�.��V,��O�?M������,Q��z@�F�ք���|͚q5����u��o���9�Af����e�V��o�R�+N�enY`�H\4���m�yߏޤ��nح�	C��hz�'���+����@��,H�kU��J|��s|H w���rݤ����XwN9��ʺ=�Ѱ��Q�8�Ԗ�T����ðp��G�zE�}a0T�ao�h���1�ȓ�I&"��Q&�a���O��=��R>�=V�ҏq��|���P���Ʝ�ߛFڀM���'C!��J�i�E��z��=~�,�Pl��Ш�WBG��GS�0�|?��Ae0~�m*u@��4��s~�GL1H��}�O���R���BtI�AJ�?�.NVW"��Z�@/��w�#��џƘ�EX�����n��ލ�%�Ko#��w�G� 	Fb�iH��D�7k4��	뎨�ºo�ژ��[4/U�NAh�Λ9��ZP\��_�-k����S����ꃠ��jQ����:p�x�����UەLQX�{婍���{���6�sVJ�=�e? g��-�]���j�,��Æ�wʥ����xm�w�eL${���|��2=�C�=��LF6%0鍢K�R�r�:^�`H��Zsz)��@��Xm��,Aҡ�p�.�� �V��y߆HlD��+���)�����d#
/L����7��&� ��0�=l�3_�}�c��t��gF�F���A@7,E���Ѻ��]�^OY�K��RU"<��$���.ۘ;������zSqK^GbNўʝ���C �M>K�n�ZL��*a��%�8���Jf�d*�л}_<���*�'�М�;[,ğiV4џ���y,Wb���d��,��v3����qF?�1�:˔��բ�����z�V���<w]��3�,��.@HU����8 �2x,�,M�������I��|h&m(ҋ}�, m�5���)��?��� R���!�f�Cw�+g�ͬ+�6�)���u��2C����&�ҽ��#�����ȋ�3!��=�_/�U�Q�?��@цS��%\f<X�V��cgyfG�����4�����V]zA�H,�(�]+�l�����%��y�/����AU�>��f����pE'�=pt.����A�d�N�B���n�\g�b�r@�s���r�K���ɶ�.E��rAm�(�t��2��t��W�!��x��e;vI�ؙ+�f��Dl��O喙33$��V�*�%�f$E�:�]�����Խ���v,��SG��=�*��u�Y8I��,�6��Zt��B�e��g�L�~շ��[��'rL�]��A�9t�8xY�T�μLE���^q���fK8SK!K��C8\�
,-��9F�L�Kc���QMtٰ.��TT��x�%�X�y�v�fsv�����!�3B)�p�xi�����D %�Sկ_��2��Vp��]�Ab�P0��M��_�y�u���	v��P#��NoY���	���{�Ul6l�����ʻ����t�p�+����wę��P�n��*��蒆d��1�_�g�{�vG.Ê���D9N�*F�"�X���sdKb�.�aO�XaT���Y6�{[�B"2�����홽��+}ʓ�ܝ���|��
�O I����ܥ&N��o���4����EIn�t8�8��&On0֬����e�+$��p��f�|箃��j�֭K޳��yK�)S# O=�~sQE�8����KBe�g������D�̉���h臦�������[W���z�a֭�����T&��bQy��i�m>n˽� �� >�:�����&���C����>�|/�������}��}ts�֡I�oˢ�+Q+�zW����6��A�D�E+k�Q�Q�av:�T���ٻG����w̲9%
Go�b=c$�,�}%ZI_��$Y�پ.����zj2��̞���f>4���X�
����Ӳ�/���$z�����U{��H	�X���~,���1��u��ȍKV�3ܰ	K֙9�4��� K̪� C�!��6�R� �;~��iP9{�Sw�LB��nf��C���L�-�n�)��L�?��'�}зk�V'�z�����8��MV\�> �O3~���SY����!�߳hw1Wg ��' ��N�M8�X-Ekva^)��ؔ���6�{9QWlX�¯�Q@��L �Ee#�d,�����[���2MLS6oo�[����;�.y-/#�&��d��i%�X#�Fr��,�Dv����Y�D*��l��T�rڮ��	��/�Ζ�д�RG���eU��I�W��G��P׮�RӠ�充�+݃�@C����+��-�9i������:ف�%]���(� ����V�Z� �~�=�U%�?@Aϸ1��ٽ��MOɬ��݂s�۰��V	H��-���V�`O��4��{A6J�sm�PeZ���7h�\>���"5�l� �����m`�jeM�f�v�VAN��(��B�H�FK_T$2@�H$�����s��!u\�rW�J}u�<˱���rJ�&��z�t�7���Qx	Ck���ɀ]-�nI�/)\�"�Q��PG�3y���ۖ�C'�Xs���W'1 ��4⇶;���q�.]J�����eMj����{X�G�s�A����7�=&�?$.��o���:��ɿg��˚���R����Tq�G����܉}����ƶgr�yP�W���.�R��+[��̸���~�WX萠7O1$Nqή�����~� =ޜfX �o#�B��{�V�C�B�S��ʄ�:v�d���������#�&���D@��ۅ+�ڠ� ]�����[�z]��I��������=te[�[�ހ��&���+���9����/D�4M]�1��u^$@�b��P��]��m|D�\xց�SyҦY��C�K�"� �:4~*?2@tG�+1�m	��NB�ur���y����5���.(��m�@��m���1�)���"KE�W�E���q��eiv��� ͮ���}��ak�4���?;��XUn"��"����L�ږŷ$ԙ�����#O�	O�;���UZ�m����MU'g	z�\-|Q~2�2GPD�0��fe@�$(�g!/�B�O�s�� �쐊 y(���%o7�srO��}l�n/7�%.�(:h\��L���x��e�? 3��((���s!A�V瓏�	�w���d�=��sT�Y��S�2PQu(����p����b]�0�nx�J�002HV�O]"�ㄳ�G�D�G삞.��n�r߀�%��jih(��3<�p�?��֙-x�crZ�4����]�B�W��Hʬ����~�d�&��?��"��ޘTS��s[::����;0Q���'������繍"d���$�b=���ũ�˧c?��ũ_K�b�,��v:cpBw�Ŏ�_���g��߉����;m�Õ�GR��o�O�,sh& v���3���Ư\3愼/(VL����JPOrv/F�e*-j{Yl��E���~4g�sx`��HTyto�.���ͽ6��3�^��Ĥ*��%�阄��яD56�`.�GSbŪw\ǔܤ!�"�xJ�S���b�.+.���8�����F� M�;�հ<<��I���h�1��.��eB�(����E\�=��E�����^]���ɮ����K,L�4a�R��Q�9����)B�=qb�bZY������o�L�?�S�3`��`�Ȑ��Yi��ԃ���.eTS����e�L���b�4�Y��ٿ$)]�����8E?�1�^�ne���ݽ��\4C���:mE��sOs�`�U�R2�S�Dkb.gE��uD�V4�:k)zr���nG�Ժ�j1��`
�˙�>�UɸI�ޕ׀�}���"���� ��B�2�Y4�j|\��x<�bO`���q�J�n�WŞ�^8�q#܌�eV��������v` 2IR;��պ��f��:��=�:c�jq�Voi18��73�!~������U�Y�E:����k��8R܅��?��c0�sR�L�豪�=���Z3L`š���ь���HDv���a�HҊ�AȰ�U&A��X��Z`����pxDV�$��{Ӱ$�<8�o�|���u�� c�K妩5VJ�]
�ݛ�)���cC��)u��r�{:攼�<����%���ש�Ң٤k�Q�
-�ԓ�{&��wg��LI����s�C��2?�����0&��v�4a|�k�Ͷ�+5>t����d�?���eG�N3�IM7�)j��~��&9���
~Yuq��K�
�}j! P��}Uʩ�mB�</��D���f" �M�C��:�ɣ���l������R&��JA�d��{vK��@!��E��8�w�C��,�\"���i��?e�����(O4�6KC��tF��+`n���,QYJ�$H'yѣ$6��Mi��>��_>�>��QaG	���p�3��mѸ���vaT���U��6
g�|Ȑ��6��8��M�����J�y��DM.a���Ϭ˳���l��z�*Š�����n"\��Yq�;΢�k�~�<d������$/}���DeNFAѢ�ʓ����-�%�;�㊯I� �C,Á�(<�l�~�ϗ��kn�����f^&W@��ڴ�엘�Xt�����8�o�sV�+Ec��̯��`�L`�j,������4��?�7�w��!��*�+J_·�)�C�*<�<i���8�z2�Wx��57��M�M{��]��a�ʹ�v02nZ�T[��e�u��F�β�ϛ�gF��À�ci֊�*C��?!�V�L9~�J���^�Y����f�W���]]m��c�L���u��ſ�g�d��$N;�L�5�?C��`��ѐV8Xa�F"��h�2�֓�c#���h�sb)��)t�1w=��r�5/f5-:�F���ua�%O��j6�`i�#��ۊYl���k���s
��"%��L�`PI����5�l�ɚ�z�$��>�T�Q��i@&Zm|%,�\T*|�eU�� �����,>�n�@~ObL���ӼU���C��Q���K�C��p򹝧p=�-�'��uao���l�4�Te�:i{�
_�j���Јxzh�c{ע���m%�q���vgiT*�Y��5���%�A�����7@�{��XF���7߱����qu�]��Un�_>[{E�i=_t=u�8g����m�����"d��%>�<d;�(�"U�Z!�X2���T��#5�N���dBL6�8���:�$��R@��L{���\2�����N �6c�23+�h����u,Y���l�`���oW�;�Ԙ�zbl(~�l��ﻅ�r9����������~�����$U�3d�����C ��H1"�c�l�d��A��8�<k �Fи%��Xv���H�Z�wT��)قz��ʤ}B u*$�t�'�𚷗���<�+�I��Ęp�B�;�^9��>�֝	6?�08_�S̈@�S�M��M�Ih��	/�,d14��J�u�0d|
�7��%a�~?�K�5$ٓ1=�5O��4�OQ��@�ʠJO������NǂM߳�+10�����e�������/�P�`�-�?{�*�J8}}�L	Q�̢l�#��%%P}�ld�ޝ]ԜN�F��Mߜ<�J�l̆8e��=���r�;eDW�Τ� Kq͉�W�=H��z5櫳_\~�!)r(,��� �ͯ%���Ղ�.��}Gc_<[���8��-8���ߩ_��O!��p�����e.��K#MxSkS'��÷ؾ�)�a&�e���2|��-z �f�p��0ܝO@K3���cPl	���Ž���<�x�6F�Sυ(���>�]GƂ��0O���嗜c@2"@.�3���_0�u���*?!]N̈́��U�^��,�K�'�7��r*�C{���IKs*u��Ύ��0������q=ဃ��Cb�Ik�[ɖ#�N�.s�r̿�G�S�AF9qg��IU��M}y��Jt�0�/Au��9}UN/�uN ���v�Fㄥ��iy��jZꅞI�:%��S�1��L�z���?:Bm�-��e�G�ư%�.`{��؉��J��;�"C�*o @]v��r��-�e;$�����rA�[���	"���|$X\�5��g3:k�mC1�a��x:�Dp�xl����J�	�`Ɏ4��*�	�O��9��w�qB��.}�cB�ј/?�ܿ̚�[&�&)��5�X�y�D�� �Q��XǷS��Eر���sX<�O���B"���d��FU�:N�4���[���R[�ȱs�a[3t��xD�g�w�>� ����X�Q	&��5ڗ�kjCdֺ8@J�!�2i7�ί�Sr�L�<��[U�w��I�����̒V[8�"�g�(�sk4:w�c�jmx�ؤ��ac��$]>'|��v�#�~[n!]R�`��,�q�of[����)����h�kCXg��
��Hbx�1��З�J�`Go{y3��<#��g��IT��ⱶm�	�`&:���XW��H�z��I�o�`g����hSQ�cꦓzM޳�Z�\�wGd̑��@��<U��TQe���@6}�JW�]vy6���@��]�`����\=�Z@7���Zf�ʅ&���� 8�w�����[�k�Rq�þv�N�w9u��;D{���b�&�ȭH�]�Ăd�@#��'�>���۝��E�_�\A]�JÂ��>wW�������'<��Kݧ�����7����7~J��)�T�h��(��1��{B�~�Bma�wk��o���'y������AbLue��,��fc,����N�W9��Bh���5�-������T�o_�����J�+h��,��+��S�#œ:��|�F�	]��+@ۢX�����MO��_�������_�8�&��ـ&��^���j�!��Q-���Z-b�«:Ȥ�v;u#�f��U���/!�Ž��,Ȕ�}A�n�q�_L6HV��|պ�E�a�A+{���6����gӤ�L^9���'I&����n�46`xR2կY�r�d��"�4��6�����}���_z
��=�_�1�r8��e&ä�${��6X-��M��2)$*�V0t�RU�nʲ��#:V4<��:
i�(u�*Tp��*�[��dH�����r\�gלYϰ�x	��s�1K] !#-�f���"t&[�	�!����>�*�Ԕ[�J���p�M�,�O`�ұ��됄PV�PiM��iԉ�sȼ��E�b�+8H�i�b��1k��]k����A}�D�/P,�9��3�ކ	f��1'3��K>7`L��?�n�u� �,�x����`݉!ȕW��� ]�gƎ��#�~��,W����W�<���G{��Şs����thD�Y���L��]��E�rt �X���R����⦓�y�㓅V!D��j���0��0�X�Lp���mU�8�*N�����3�#��g׹�dT���^Gh$�g��J�h;3f��z����~�i�
�w����}6�R���[÷n?d�ɓd���nB�ۭ�h���>Ux�4n��{�����aWp�GLV�D{���$�3g��
��"�[-F�\�B"u�P��u�s~(�b�>��2bʘ^������u�7+[E�[-�Å��j�|ێ~xA��G�3�	���61��A�o]!Kn������Ӡ���~E��!�.ϏY ��6B��,hv$����5������Μ|T�h3������ >Y}�t������3T�_�-6�e�{y�(���0ѽ�HПP��C
94��<���
�Σ��w�C�	�pFor�Q�B����vى�����I�ɯ�4�}�pA�(��>��2/���:�b$���_��q$T�Q�wԪ��Y�Y2�Tl5,�zY�k��5�p5<� В4����icӁ䘛�Ȉ���&Ũ������9�i�
V:�վ��|c�t�� mCK�t�/�V��zg�r���Қ�n�u]��m���;k;[����4����<N*%V-f��5����/�ӹ'�!�-���C�&�>��,����M��^���] �����t#�ׯ����.�X����i "΁�4��uG��*<o"%[G�9l,_Vڐl>KK<��߼���q�{4ݹ����M]�����i�
Υ��H�v3I��Lu3���)�ף4S��1+�W	3�qх�����v	�}&�M2����ӟs�Ő��(�aZq�+�gi���E�E{�`��F��K�zƧ�p�qP �R��K�@�p�$ [�K5H8'�r\�]��%7�,nR½ՠ�q�����!eK4*�n�h)y�S�����������vAE9;z��9�˝���u^"R�s�� b� ���+v�x9��F�J�{��@��ͽ�i*EjC�K�f}B�F�*r�Mg5�A�էP��(#@�K�L�ы�X�����H�����#OQ[ҫI:	��!�+&�9Ǝi��V�tt�۴Nx��@L�k*��t�v�Gj���k#m%L��@M�}�'l�����M��qa���9s©�s�b�Z^=&*to�u�j�zuo��l]�YHo5�0�05't���.Hi�ټ�ʈ�E�Cy�x#5�y;�kt����˴:DS��~�eCW" ��R]�{��&>���D^f&���J0%!�˄��t��'��Q%P��g�y9���x�jz�����>�����5ҏ1���'��H��S��zWv&����!W1���aݳ��؎�����q|ä}�j�ZC_��@���[�|X�A$E~���r�L�R�d%�ma��<���k�;T��������r[��7L����t�=��e��⚜���CҕL�^n:�����
����X��̩ͨ'x�@���t�\�)���;���{1�������ni9��l�ô�dģ-�7�����kc��VA7�ũy����n[��*_�3��Ku�3��m��-�o!Tf�uEC�?�X8̹�O��J͠?��� w� �^�(D���/��xmt^�� �Ps7:�G�h+�N�K��B(�H@�8%׺�58�?��{��H�a�.���#��tW�����̆�Rf�`�@�bf�J'�Qp]գ���s</n����1� ��KRX�fk�,eo/��t�$p����эjD}ZyĠ3�����m���Ի��c߲-����k#Q�!�p���e�"馄h���{��W%ݵ�gJ��.2��I��+a�S�� �sH�ٰlt��:�e5Z��b`�S6dx�~�uNKyg-Gw�ح�a~�E.��8)�Le2#$���
d���z�(i����	5���p��K"��r"p�Cob����Y�=x�f_��у�e@$k�c�0ү��.�9�b���ٸ�aΑX�m�Ao��`�ݵ����m<�s���eJ��H7�j`?�v�>

-�	��Od��q�n8��t�`���dzÔ���򌬷�b&�j��o��Z�(�g*�ŹX�{�؞w,Q�l��Ԟ1>H2`�]�\xq��M0`��ܚ��t���G�]�Q����e�j"D@��$��\�u�c�3�4�̗����V�*��>��#��b���v۽Z_�e�r�L'9*�W1�z�ٵ�jf��o�_������p�i�����u3Z-�epK  ���C�>�7��M������b ��Xk0�UˬS�Jz�5ZTz��~[����΢��n����-���Vu��]Ju�S���������!Gn2�"3��6���)�<^����������s��3�C>C_ʫL� ߎ6���8�;m��6,��%ں/~�
<y$*\�MYㄭW�M�*@�{���Y�y�D�>�Af���4�*��������{�ʈN?����#X�bc���r#�4>��;��ef���|��DM� 9Z����	��|����C6E�H�Z�T�L(+��菹c�!{����?c�������j�a6�z5�EwĆI,��E��L�}Փ��	���wVn�7�@nz�a�&�� i;���ӥW�"־��>[ ���m�++ �C.-�����c�W�$�����f���ƛb;���>�O�2O.ʵy��I���E��H�RO���I�l��ܨq׉�ǥ���p�C����;/��E4�jki	��3;�Df�(Q)��z�$0��h���ˉ�.M�b-�����a�l��;������J���/���yp��2�yβ�O�Dt1�WC�����Xk2�\���o��
�Z�J�	O�[L��F�e�v���ok�DɊ]�3�5WdpJ�a�t��+���>��/z8��������n�]��#I�JE��k�����h�-��ڠ����)K�s#���SC�s|��ǈw�ʌ�)'�N�D&D��'+���� ����T|��TR��RY0�k�����-�����z���F�M����]P�,���\�2 ��M��[BL��H*���۪_:���U����m�$��v��2�B쯬zy݀�^�3:�K`3���7�;�~Y��jv��{hY�9����.u���!�8ܟT}��^��N)I����v<��h��\<� �>47�%D�	�n~
����Mʜ���p�h�x�I|A޶/��ȗ���SY��j�@ ��V�������)��n ��R�2;4Ջ�f_�Y���
b"�)0.8��6��&��@�R�ل��d^����I������U�@+ &�왽�E�r� �ՔdB�Y8kpx_7�S=�D�B鎤�����+�6�l�	�7߬=�h��f.C>�����NL�ye��p|"�_�p�_U�j�{apd���g��+{�;]^�G�j��&�n�F7 �Ee�2�=(��UX�_���gG�g�t�~;z �lfT�� a����c��s���@l�����d�R�V𦅐������>x����đ}؞�f 1Dw��3{���C8��?�a�Vj��cIy쮻�0�W�}�����fٶ�ZHF�BX�D�S���rPK8�v"
q��[��cy	�T�_f�����}�ةX~�d���F��������e�p.�����b�F������I�e"h ��vK��Zd�H��7�ԙ$O$
��U��9�fCL�0���S�a����s7�wp����-+����j�$q#��k����u2z�d\�\kZ��\"�(T���p�f{�Rzە����c�x�'��17��/W��z�� N;���[ɫ��pu��� �^��a�ů;�{�K8Z���ֆb0;(��j��}\��!?��p3�-��<�f��@�l9_��+豓gx�)��9v�+D�
`:�r�ܐ��F�]02q������?�o��;�śx�r	��X�T�p�χ�Qk�h�H���z��$+,�gZ��0�ܜ�PbΓ?!ꅨt.Q�e�k!mб��OK0e��zF�+�Y�4���*�����@��ݴw./�Wd�3���.��-���A[�$�f���|�/����F�W�'����F[�e	����0U"r�T�ߩ�>{��#o�[P6Z!��&��t�3>�[ &�5����@�B��i��{���{���V��z �6�t��8N��|�f+��"�����R-��[s���?	Z����`�Eg1%�ev��$��v3������DhݞKs�"oOҠ�L�5;D���:1l/~?����g�T��$�mXTTGvN.jh�*�OV���@yv�7j�oV�`7�w�v�5��3-���+���@�bqB�Ii��ٿ�5?��8���tf��y��v:�������]�1a=2C��"�����O�ˉ �oy�G�J�?E���'z� �H�pp:#�Ȓ�1�E�w���y�0 X����Q��<'%jI��s�.�f��`��g�Vh��ro�O����]�e�$��|[��VT��nQ�@X�ˏ�t��t(k�c�ʤ�KiW8%���#7lhNY�Hx�:vxn�2.������f/��u9}mHEK�����o�-��[�����ĝ�1�y�y����_�ܱ�e��
E������Q=�[&W�r(+��p�;I����O������Dm-�hxyVb�癵��rm�?�-��C<�i�$�$�CPY�"����W�v�dKB�H%�'�X��;�'Y�{F6k�J9h������_s�
!|>�!�5M�E�?��ȣР�D�tb`�V�k���i��ß���fl� &�l�o5֖u��z��e�K	���:=�����P��۽?,��3U���d������pK|�����y���������Eo|<��`���v��b������1j�'MR��'�,�R�"	!;͚Fk^	2 ���}Kw�*E���W�y0N�$�'-�|�IO�H���-�|Lܚ~Ć����^�P���2�~�}<y��bF"6��r��78(�Y�R�1��ÙAJ1j�p=9�9�\fm�e>�AD�'x�>E���ӫ��i�Bn0}�W����Ķ��Bo�U6�=Ҵ:d���䴠���H����~6z�du�A�ߛJ��+2�q�1	.�Y��P9�e��%�"�z�Ҋ���9PH�b�y5�9r���$r�~{��Zj�{����-6{�l���j�H�^�A�R��1`29�+8�=��)n�x1`���C7<x����s@հ�X����.���8\���A�2��0Ԙ�x��Pۘ��%�B�~p[A��$	�����|�ޫ�_�#�֢TO�ǯğ_'�h%9�*��[�
���;���ۈ<-w���`��8U(���DŤ1����t�4`�"�����'ɚf`��K��������/es�\v��fw��2(�q]�t�p�#���JE0�^�V]�g@����=��H�/���6g�kn��^�״ͻ�$�9��x�P_6R���z�,���G�2/�n���^��e�_­����__������Ps�Oa�I�w������9/�� �ár���|"�ѷ.���$ё(�R��]JZ����W.��S�
�@�[kv�n�"*�Ҽ��~9RW�����#�뒏�>��h@H4g�H��Y�M���ǁX���;��*�y��ـ�@��k�Z�Ԁ���\��^�I0���	��6@�H$�t�/)���.%2h��z3I��^Q�4I�׼ǝ� �),���`�(T�_�8�_���{ɓ2�O"�����XW�g���+)ͼ-ww�UG)��߹D�ɕ���b�3����/��E����]]o�/����f�	ňE[Z[A���i�ċ�E��+��x�V����]AT�����^KtB�R�8��b�$<ѐ�V/;�YՕ��LK*u�� e���ky�%���R�.�
�Ak߇�KߴJ�:�5�5�C/Tut3��wL��"��:�_��A�^���c�H��
�B�����uwX����|��8�zY:�4�!n�ݥ������2WW`:u��-���<��J�a �!!�����5��ߔ�dŎh9
�|Ҟ�R��e��z_�e((}����ƭ���ܠ�b���+ +6�i�`[L���z5y!�b ��J=gU��zֱk	�y}	���YaV��jp����^�mD��_��Mׄ�r&d-*��9�(u
�Nč���|T)m5s����$5����㿌G�
�[�za)��O����NҺb��zT�K�u�a��a�4O�����)B�3�Ģb�v�u��m#\�(2CIBz��:I��i�n�r�k:0�eLׯ�'���ט��!X���j^G}�V��4���#����P��rfP%��Rla�j8�Z�K\�@8�s	NWT��2lP&�f4��NF،�h�j�=�H"�Ʉo�k	)Q�4�c�Xc�W�e�:G��@��W�<{R�m��(<xDs��B���k����]��5�yOҏ���/ޅ�i����G�н�Щ�ճ��E/�NG2淎`��h�2���:���+���-z� kz�~�ڏ������yeS��^� �y9CAhY�d�]YRke�_��ڲ����?]�<S�X�`��$e��u��ݿX��Y���"��F�`F"�/��M�K�^d���{�hm�j�k����櫏5*���v=Hj�����x�(#S��z"�>$A���J�~��$�<3��w��y5��%P�5���f"�#�_����e�r�������K����*��~P�?α갉�<�[�"��_.oF`D�I��Ђ�O]�w�rO���ڍ��:�J�B�V��pU�/��D����0�<�Y`;��)bISUkc��?K�Da��5�z��W��x(� P����H
(,4]��ØFC7�-�zGh���-C���x����#4�-v_M�["�{���*�񜾚:d�$�*�Q=�?ĩ��+�v�������T�2��<��_�͛P�0i�^��?D�t:\��!�%�Z	�M

V���һ|�cc�4�������t���%�c@l#d\nY��݈�o^�8ѳٕg)����t:�:ׄ�c�Y<b�w�
�GgT����Em�A�{�E�3���WC!��O����nP�u���  ��: � �w���?7����/����'��{ä�(Z�i��ᜬ�־}
:LG�~j�|m������4���bI�����^�~��Pʠ�|�2����Q�8x�d��`VN{�,5]��ni)�]��G����Z����i��oY\�㼃�8� ��8"U\~��Ǹ����m+ R�/��[��_�ڔ��_��L.f�ߤE�j�	ɞA�l��.")0D�_R9��VOD�z����@��A�����Zz�C�����BN�sr���8<W%+&(2���s%�ܺ�Ҫ����l�ϱ}6z��1t��c]J��(��ߗN]�%�KP"!'�o�C��#��0��2ߴg�|�X��.�r��̻����"��i��/W�L
(�[' �tV���KUT������Y� ������y�i3�lV�T������r�n�1�yIU���O�(q���ߟ�kR�,�"鱎T��w�HN���2�ď�C��@t��9�P���5���c� !ڃ��c�:v{������H�#hn�Kܵ�����i�Ό���+�
�_������1���p�����2�-�"�jnS(W�	�~>#���d9�l�d���=`_���|Q�6�Ӵnd�T��fx'䳊]���vN�4�<\����A���{4���˂�L��$]��9;e�Oa<�;˭2ҹ����8v��e�hl�#�{l�?�P[��������zt�м}R��y�%��;q[h./1�	��2�u_��/�UJF�33gKUFbVwbU��eY�êו��C%@�E�)��������ɽ+��k��B^"��M�8'�e�\q.	<4R&�`��n�/b%�1�z�lO�h�s���$�RY�'���Im�Gf��W��b g&���h�����T�����	N�IC�i�5h��Z� |
{�g^K��p�C��1�4��Íct0'f�7���l�RO�Q��L�W`��.fG_׮2��Џ+�Û��v<�:��ƻ&�f��@9���&�i
�pⱏ��+�;dA��"�+U���ov+||�c�u�1�:�ț~��ºYr�O��`u���Q�;��&5�a���p��L�������8��K אy�:9fW��8��E6��U�@K��i����[Wl�%��=(\�4r�{Iꊃ�"çt(�{�>��1z��[%����0�&h3�HЩ�.'"<�O��AfQ�.�]R9A�N��)����H�\-�,2w�^������C��>7����4��=��Q�>�_`�lytƙ��~�<��
����lt��Q��"��"�u�_��;P��L�r�5��@�oi�ոp�Ha;J�F�n�8�I��0��ؒ�&G<�B$UҴpk>��d+
���d�]�ٷ�����, �����һ�>ZO���@�h�C�|?l�����Ne�2</v��ݷR^;*+����x�6c���5�ɫ�pʱ��� _��ֵ�H�,���Ƣ��`!�c���?J�����}3`(H*����8̉�d`�`X!�Sp�7d)@�E�-v�q��ͬ˻p�vjkf(8�:.�_�&�x��'ٷ<ty�W0�3S��]��p.G9p�k���r�������9Yn�a�Rj�i��3�XE������T�o0�߱��Ο%,�[�����W$���[z5W,%~����3�_39ae^7�{׹�<B��?&,��|�l*%�,|����J�]��M���E(O�n��dIMv���&�,{e��ڞp	�۝u���0�A�ۂ�!؋��aN~P^�2��0o
���j�8a�\V���t�$/�-M��X�T�ym�jj�8to�"X�n��
��ص���rVS5�m��GX�f�QĻ����s�dG���H���g`0?O��K�Ų���xP�Xb��r��W�C�\D>t��fh��'7Q��]���`ܽR�W�y���ߵ���󖡝g|��|G�*Z8�k���IJ�g����J�U$�<��	"�`r-���?�x��+8�pCl��&/�JE �~���9y�W�9�m��p3�ב'���a:��8+d���<��g4�:[�'f�?��h�*�3&���{~�P0�*��]���J X��@i��*�T�}#!�Ӏ�a5����t:I��d�Ɖa:�*�0FX+w���n=P�҅�`(
�?���g���+B�����6. l�1�OEln<�BN�eʜ�/,A����WX�pZ�P��&&�yY���ꃴ`�&]�@rǲ���
�EE�w�^2�����znT���#ļo3|K�o�b����Q����戄J=e0��;'5� 2h�:���|%��Z;�9��,�<���Qd��F���&���f�Y�p��BÒΛ����-k��ú�\hΆ���r�{�em<)o8�{1:ߗ*V � ���߸ГW׷�L�V}:DRK�u� H<�;�Q��f�*a��v�:Z"��὇��������T�	�hUpf��@,cR��k�����  c��9�w�6�Qg��|�0��H�D�y��ƞޖ�s&Ǿͅ;Y��ƻ��0�w� OG��.��$~Ҹ%q/�Ê5��0]溑�)D�S��cH�R�-<�$��]��YT��]��%�l$-7H���8�?��Q<gܓ��r�	���x�-�����!�nJ]n��ȥ��B��M��@j�;���'�Ń�u�����# a
¼M���=�@k�{ۆ7��G�ހ�93��y�_��2���m�,|R���\F�*W���oOX��A�:�s`����/�T���t̍�<̩}�Qi����<?'4�'���z��3�ydy�{u����H=����7����M���,BT���3�|s	�t߶�)V���=����)��{����Fh��������F��(0���P�V	�Sxw~��3p�A;�2�e-ŕ��K�&��?�4� ������!���+&��0{�,��I�[!�Fqy��S�G?XA�86`�~�$�Y�� ����4c2�+}}��;��g�|��b5` �	�k��:�wc��'�'�U1O#��{��T���W�\\���A� *u3�����le�ҕdw��fm��pڟ��
3�$�jH�ޮy$�v)wH��M�f�,�y;����Q�벽�r�ϳ�-����@��h�'�5~��L��@��Yr�R�Ғ��E�&f��9�An��n�x�o�nF���#�L2xQD<fy"�Q��@&"9$c3#��c�w9:/s$�#acn}c�Βt�g'ɣ.�5��S@��zM�p�J�M����&Zݵ��$Yp��|�K��Co��
�c� ��Ԫ�#�7s�{�daz�w]dˈ���iٴ�h�h��	�K��c�֑3h��#|b@!
����"�+�_��/Χ4M�V�<U��V;�~w�,�j��a���G����w�~2q�dn#Kb��d9���!2J��ԇ~� �F�D����5�2K�R%x����+�_�>,������/��5(�׷ȯb����6Δ	}k-��Ad2"D��k��Y��L��=!�,����,$���ɀjLT	�0�` �lx��`���Ζ�v��	9i�D�R��>���rOqԊ7STפ�4mI?�Z��"���-VU좴#gT��Ӵ�`߲������_��jx8EU��crŐyF�Zs;8͟hA��ƹ�X�v���9�s���7�<�����������ٹ�]��:w�u���~�ؑo�'h�\��g���Xl!����|Ֆ��^��g�?�VO����zMH��X���mY_e�� ���I��q���~�+ 	�",3����8˨���p�裆�Iހ���
=GV���}�M� ���E���aC�p�:�+� ����Y���L����ٰ�7�������+_]�_��� .�hDduė�v�[�ۜ�|�j�VL��#=��)͈���i��;�����FԴ ����$�)��.{���ҩ:��R��p�tv� �������T��S�:>����ih���J7#t�}m�,��G�D(˅�&�RXL2B^5�b�,cu?���m�G�z���ebȗ?ԍ855�_�������������E0_ԩ(:J�ga���(�>A���U{�E�9nF"�1��3*�T?X��x�v�(}a+�r,���J �2Fc@B�B1��&��Ɵ�n[7�#������}MG7�w�q��XA�24��k�r���0]��m$͕ѯ�O�򹠼��,�$8�x����h�j<��-Ay�QgV������~ҧ�B'���&�qSEQ~���͌#/��D��-��6NF��B�d2�O��&�]7�.gb�@�U,��G(-�)��MB6�YAW$NyK�c=t�į���4�ѳN�����Y'-T�m��
�ZN�e���hqvaLE.o?K"�)7�U�.��9��K;��wΛ�sW�6���M����L����U3Z�jEס)U�FaO��6�>1�7�M�J)�z�0��R+�q�ui�̛��Dhd�"��|W�`��e�%r�9Z���d����N^ɉ���<.�D�� ��:�W�j���eLC!��RB(~Ь������2��I�!?�e��	l6L;A"JQ�p�����_�d*��I�VYyk�|�t^��jK�q�y�*n\��{�R����v��A��S�K�� e�:��R���5
��:�#_,�;?�Y+�34�]��\�K�T��Az�	,2�d�F���!�v�'�|ns4��[��it���if�=�\�-82��=T��X�8)&PW�xI�	W	R����NИҸq%��v���T�˃��w3*��15��H��,pX�����Rm��x��(>�fM��+op�ʱ�3kfE[�n�3�hu��ja��_j��e���rމs���c����Š�,�B�Ofژ);nc-��U��I_��2r��6���N�h�t�|^fᒨx;|��.W�FX3���h�evl��k�<V iO�x��ns]?e�@BQ.�  x��ƕ��0!�X%��@ݫ��x{3i��Y^�wS� �I�"����L�W�ׁx�O	e'|��I�*����N�)�d&����8�9_.����D��I�+ �H+��;:�it$��Rψۤ�B�Qŵ��>S�<7]�!C��?��Oۜ&9�s�\�5~j(icI]E|���d�ɩ�'dP���C�Tɂi�d����SRw�ޗ�`��q�/e�+w�O�� ��	��[G��%�vF� �m�;�p��YU�~u��֏<d���%sp�TA-4�\h}���H�C�~|t������X�Ť����Է$�<:M{μ�Ql����Xk��U����;���G�q E��T_�/T7�&
�r�6��m��)C�> [I�*8�a�g��x�B9�%?+��Q ����S�[����{z?�oj؀	╺���9畿�c�c����Kh@�iЏE�;2E���5��.@ߓL�>�2�r��O#����M�9.	=>3U�U=��?j2�,и��u$��U�5�U(���e�O���t��7é,�W�f	+5���Mh��T�۹{V�̓��k���"8�����{uk-
���TK�]\�� ���s������|k��A[O�XH��lB#��\ �DTօ�:�\�7א�uiQ�8G22��������A~@P�a��(�D��)�.vl���7P�s��y���:L�M;�ZA�G�4���u���y���I�(�M�F�ܝ'�ͪ=s���v8L�[�Ѹi�~E��:.��:�Iq�N�I��1�V99CM��
�["�����e��U~/q-��v>�%�zO} �u!_L�Qa��[����w��UѬC�Dg~E���G��L�,�,>u锹� ��Ul�P��a���q��M�>�ɷ�M��C�hۛ��S�bAG��d�S�z�t�:�[��u�x3!�P@�}VpY;�B#���rY�cwA�kݢ�`��sڒ�*��%�0���4���MhLq_`���� ],�W�>�b���z��,lVc�LG��z˫|֣�L��l�+ھ:Ws0�،�1o.O���̥9i�&x�C��?�--go~#���rNnV��.����9�u�v,�2*��Ϥ� ����_��:���@�,���l�P m%F�cw� TgK��<A�L�.�N�d4P/��?�1��J0�w��z�Tj�8�r=�FO�%JP���x`XF�x�~�a^Mj�����x��Z��\]�!܁�5�EBJ�����S�P�;ee�P"�wb{1�O�n���&��B�m$e��06t�]���4.,��̍�>W�$��*-.�k�:�O��B2�N/!:f�Z�Sϻ�0�E���u-�Q{a�E!x�&�tڗK��u?��B�����HN8ç^�7r�s�P��q���Z )�s�f0	�����6o�5�&k�Z���.��TZ�e^�@b��ך|���4F~�rU����J��?#�4���㟶X���A:�w��4@�7h]��Q�	om�me�J���a�v>���)a�h����V�oy����;��\N�xh���V��+�� 7{PY-���H][��Ƚ�ed�nѓC��$��Rf��$P{7�O�^@u��sm�%9¸��Ⱦ=UBą���^��%tZ4&�u����T��&8���:��B�/�������������@?�O-�����d�ٱw��HS�־��g&5T�7�p��!�QB�O÷�\��EЬ�~�����u��P�7�U坊��J�z�R���7����W]�k��:!�^��䴦���k��c3��l���t�t��X��춛�
L<���lP%h���\־$dc�́���/��L$;叢s�*��>�nUo�h�����a}�佻 ��KEt'�I`B�����M<�y�� @a�BX��K遷��z����I��5.�3~_>h�d3�襦ZE�< O��T��*�>��!��q��V8[�Сz�`()o+\����/�輓�)V|9�%��>$�Gi?�G`�Z/�A�!�
T���2��K���Od��g_�Ɉb���������pBĄ �z�Y���R��>���_� ����;�FQȻ�^B�z�zU�F�O�qAb����]�*�y��7��;���ռ�l��uTT5��z��l�~9��2 #M��\�5t�oz���ŒKV��K-}��E���11��آ�*���¬�V>�Pl�ߙ��EP�0�ڇ�/�'�{}�T�2&j���v�\a��ퟢ��K����d)&����hC8AG�}?��D9�.��Ŧ2gp0cAXs�S�O}<=gM7�&ؤ�z�d��Oe�҂��>e��QxSY�Z��@
���ƀ �~�D1�\��.:��yh�ȱTY��o@�`���_{���{�#�Bz�,	�7����ܼ��Î���9kֽ�"&���Ϛ�N�H����=�k-�R)��M����3�0��ȩ�Y؂�	#�ޏ�\=f;�����w)��D�;?@G��<�Q������#����ϖ
!=�Lf �Z$����Z&kgU(��X�ZC|�N_�}�=	6���M����H�f�EAv5��_w�P|Xċѓ8z�ޖ �T!���:�8F-������E@rZ���;U��q��7$��ٓpxn�&Jk���O�(=�U��?��ٯOF%���'�o����t��P�|��a�i�� ��]���W̻Y�Y���G(~���!*��֗>�d0Ƽmd[l� �)�@���i���.-<�;� �UP)"�.f<T�^�'����	��7ڔ���D�B�0l:IIcD�u#g`Z���5~����ڱ�u��';���$XMlMi�$8��UW\ÈL���N'�P��V���}��/��d:�{�*�#�[ϔ��]�<|
�&I�ʯ^XB������A�9���~�Z�X61IC��?�N&�O���q����&�ɛ�9��v
�U�`
���^���j�����h��k�a Dу{Io�}���"F﫹���|�|�1�v1�C^S������^t�Q���'o&�IIl��+�t�`�<�B[�Cb����ЫdkU�~{*�p�X�����X�_,�R�}�'�7J�H��R��4�hra8�
�w�䘳�Ѕ��J*�vi�PI��=�mQp�����F�W�`LŜ�<����ȬK��$W��:3�U�Z����(Z�[N��JDy{;��Y&�"V���ǟM��,�X��&������e��)G�B��K�%cD&�hI��&G�s�3��P��߬��B�X��%�r�dLd"\{�ՀR�ױG��b�?�(�T�9�{�^�����.pi�०_����EQ�'?��x�
[�6���s|rH��� kN2f$�f~��r�D�l��>���v���V��u���>v�$���	r�/@;�z�Q)��Y�� ,�i��+p���lӚn��1�b����|��*;�Y�q�"���?��0��q�-�F��z���	��硦?��~*1�rI�P9��H+qw	��^��Cv*�<d�R{%�B��OA
��f�S���\��-{��]#	��b�#
�K�RFZ�UU��f�/����w�|b�����\Xk��6j	Ã	����en.�^�"*�����@_�����r�:ޒu/΁�؂٣w����t��|U:i8����	W(~LI䣼-���ѵQ��M���йX����A��D�et�1ܴZ3Z�Z�8Q���ڼ
�s6������2$�W�H�?�̮V�o`)-��f'/=�?`�u�ohP�V�U��<�O��S_�[�r��{�d��;��ӿj4%8��µ^�C$_�n�p����{ΰy%l�I{���Ҁ����.��?ц��G�_+��X�msm!��)F�
��߳@�=׬�M"_�4�EC�W�r.�i<)a������%���#���H�P}ǯ6�c���a�P@��t`�UzԕG�;��G)~H�RO[�!�����T�0y�~�#�íY�ؕ���9lO����&�F&����0��	�B���=�F�2[>9=�ˬ�bQ���j�������4a�������f]��J�K�V5�Q�֠X^-H���MbYٔ*%ظ��P#i�T���\�����A�{��j���%���A��Ƕ�)A�+�����Wș|�R� x����3ڍ�*t��J�;-���% �rl�ZKW�E���c��ε/p��kIL�4P~xa���=�)os۩��\��BůG��>�&���nmj�9�+Z�:��(���0D�8p� ��s�{��;3g��8��/lC�.�;	��+j������I��%Q���8����?�]����@�wv��Sw[s7-5q�lx�����w��2�J��ˎj����q�|�G���E �'1Hw�R�f�V�9a����O��X/&��-W&O�#�jh��S�r;��ѝp�o�ݧ��ޞ2��&�;
@���{�7E��@��������N�0�� �a|�oOS8����1`:��e!AzO��.w���t6�b�J:F}�,��u�M1R��9�W���|;�-�^�u��� ޡo~�[��qm��K��cط��RrK�PyIQ�c�I�#�Gl�ԑ�f��p���ʇ1$0}�	�M�.v�B��]7����Ed��d�1�a9�7.���U�j�P���}�}��z���G�貮��L�'�pLI֬k��d�ٓ�Ϊ0�OOPs��o�z٭�~ �JiM\W��:�ؾ�4@�n�J�*Z3dD�6��9hgw�+������梩 2p�R��F�9�yי�B� _�@g����i� ~:�����V���H�9ԏa�p���m^SrD H׏Fv��s��^্�s��<X�b��o�g?}f�L���u���}�[j�9$	�㴩�K�YJD9��݆�u��y�,x� �>��6�a\}�Zc����b�$�^�H�2D���kdؗEؖ�V��n3�3]P���#b,U�0�R��-#R��cCM���{k$:�%�����е)m"�h�4t��n�P}2�z��.i�aJm�D�Ts�i/+��eh"�v���&}���87�u��~���
� �p����C���,�$I���I��H���BpBN�dUm��i˱f�����1�J�:�J	B~�,E�C����<�?=U��W��m�nOP�5�i�d�"�F��<h$,�d���M?���8@���N`��WA�Sdӈ~ ��Jw���9����%�S^ui!��$w��ޣ�Lڱ�屟����
8��ګJV^���a�\P�\uy[{I�s�\�����>}j�Q�hx7Ӵ�V����9`�ρ��-qܧ*f���n{��XW(��G#�����_��U����C����%JGC��X=�^���k��r��/r��N�����3� �z�L����ۨi�~�)ܦ�ր��'�L��yhN��I}2d��ا�ځ�U4���o� ��N��O^��G<�G���x�8b�m�C��WL6תr	��L�zWMC�0����S��R'�����*�a@�5U��w�8wX��әF�NV�;�T\nN*�z�
��IṄ	�����{^�_����u��y��ŶK}�=f�k�GeB��C\��H����5�(2�G�k�!�����bĳ�AhÐ��w���Z1�*�#������*eWHSr!zȩ|8S�+�����o&ϥ�X�b���3�	+�h�F��Dt���Y�:W�_&�g��O��C�t�����iVw2'�FI�����k!,�H����JcB����t�U����3��Fֺ9=߶MY�
斏�[������U<�!���%M�N	!��w뙩��_���-��=:Uܝ�/���?=����ѷ���6:�dI�G�1�_�s67�\�/�n�܏�g�?�����vI��:���n�����Y�4%��8���X1��wDrJ��u=T�?��*B�Hҏ��l��������r+�ĵ�l�B�ag���n$N�'��nt��E�j~�������hfinx'�y����_оq�2�9�,��<3�etlR���1p�Ф�فӶ��o�������l9w�l�Al��vG�-��I�7��[�lnj�ʋ����3��m�`ĕ�t�՞�����7���#Q߅�+��3Ws��Of��~>��W%L���&9Hq]���������o8�
�=1�tl
�+�S��<���0���U"�78����,T�_��!���1��}?֍�Y����'>qs
�V�r��@�&9��w.Ҹw�f��X�@=���Cj�0Q�MP�(J�X|m{���+P)�]�Z�$o����)0�(��u$�Mm�y��^�Nq�U�E|Tܴ�)�APB���:0��Q
�J���ַ����k�AF��Fc��'�>Efm}UXⶮLǧU�$x���'� �FI���,&��5�]j|r�6��]��
��1��Ҏ�s�	�Z��7�c-5l6.!�#K��%-&@��r�,}��=��7z�-67�~�mb-�ͩ����;�C�=<i�@%t�c��e�>#]c8+G*2��Q�� хHH{�#�k^��C/�AIb�h�R;��}�[2e[�n]��~��z����C+|��b�AN��D!)(�eC_=j2�Mlf"њ �Ԥ�D=�j�Q��(��H����*)�+�����;{S뻀�ö�#_�܋�,+Z�.5�Ծ�<�!b[���������K������J��c(0�6?�S!ň�{xm���{�<��DQ1"Eڼ���ʍ���Zg�1�C����� j|�d��k+	A� �#�X���O۞�2��y�������(�Hn��B���Q!��]1��A��}/P��y?%O_Ev�4rW��稛�9�f�0g�R���dBTlϏ�ߓ�Wr��;��}a�u���+�03EȧԄ �9��T0=Ҟ�i���B��qȽ���k����Qe�KV����PV�a��
�I���#u/��r�t���UD��w:�ދ�;Կ�$C�_�Ɨ�}&w�Ɓ�y��������_"8G=d�#�]�K��*�3Z,ekR�B������>=9Y��{Y$a���ޒ���y�i�V/L�*�]���]�c_%�1WW,�������\g��>��/��P��%rۙP�?��p��YT�q�
 ��6�`N�Y�����b���]C����o��o^����^[�ʥ�e$���/V����^� Ű�(�X��g1�:^vU�g�ѣ���� ڲ]$��E�}R��H���hH�Y���+��K#j,���]�`�>������ѽ�J������wŧ�D�9�8�I�ҰOP�+0ETr��*�}���$Mx�L�����dJ����խ�������	CN�%BTɈ�u�ٮ��;�9j����?p�J�$9#��������lz��13���vύ�ږ/�Na�ϼ�H���mu�w�X�����㺻h�H��/�/&rt#�O}�����7�8#�Zdek���rƬ�����c
��� 
w��tc��S������>7�P3����@l�����,qEBFT±Y�o��Y�#$��9G�e�	-�2-�`	����g]����M[*��֣��=�S���(��6G����G3lb�z��%]��kѺN�/��ߠ�w��S���S42��)�(� >�:KC*�x+YZ���,�C�c�|w�l1����F Vt����9���	���� Fw�������������J�W��.׍�4�=h�7J�f�U�ܢQ�9��UM�������rF ����u��	:*}U�Q��N�	o�h*�!������si�x��i���6'���)±8��I�Xӆo�-��ʺm\Uh�d������
N�	�䦭lsF���ө%��xV� ،����U!�r�I�Jn��ל"��<��]1.�0����y�Fz�=�8sb��H0�F�GH;/�Z���bi��Ѿ�'������D��{a����l:�6ox˒�E���^�[$Ե�?:�S��Ӗ�6��Ô��Dv��8�ŕ�(����#�[M�K���)A��H�:����<<]Nu���)�ɲ6er��v�;����)`�ܞ%���s�kz���4C��c5�fyp)���g����g�1�1/��R@I�w_j�$P���QcR�k"��p���Pt��-���j��P�z@�Z�=�;�ͩ�o��t�����;c�|����\��׌��3��u|1:T����8,�"��q���8�S;Q�,�LϚ�nY�K��pu ���-��e��r��VY�Zg���?����.���ϼM�>��5Fj�,�w��:q�].��Tp� 5��&t��j-9~��r�9����wC
@Ӎ���p:�"'z�m<�~�˙���!�H��E;�Dx��s�{TiB�@�io� }�X��ؽ�h���a���Q��'��#�5cY�1~u�� �Q��S�,3V,D��8K�_�ô`��������
B��&�PrGU+юb52����v�aʰ�4����o��n��C�]�<�,R.���HB��	>��`�(!$k�I{�-f�-�E����q�oF��
��
�A`\�0��Ɍ�+^�G�Gԇ����0�|^���|��֔X�4/2ɨ�g2� ����x"�FC�2��*���?���ªc������Ŧ+QB�%�(W����+����:��E���ެ엯�AX�v�MV}
�m�M���'���<݈B����]����B��4���)����p��.E��)�L�Wq�#��8�q&���޺a�J�t(���ji��q��G׌�}�.E�p(�;���vR�~RrDx�x���W	bDm2i!�����PY4�
�GC}�\�Qv23�\�cFmś5c�A��s�����D]�,�0qs��WCJr��G$�(��
(I�#����NZ��`Ųݨ��ֹI2g�/��-�
rE7-�mE���b�c�T���nmq1�E����|U�	���!߯4���q�3kk~/J9�鿐`7�y?sI� k�Sqؑ9�B����-����V��x�jI��cT���@���o9��>bctV�y��t��í ���x��dQ��Q��+�:a���NS^�Y}�nC�Aѯ3ߩԓ@Be�<�.��]��2ЭpU�k���["ά���P��z�p��jT��V6��
H3�����4�:r���^V����j�R�H�j��7��S]�g�����W�Q��\��B��)P�6�4���pfh�`y�W�Uуz{����č%E-3X;�#�k���__yp��x��`�����1�� ��Hz�b(ڊפ���cxu"�gY�r�%���gm�:�mҒj�k]S�&��j��P�a�6ݢ�2�K�t��%�^|�Ȧ�7Y�4��}��।II7�sGx́�AA��d��K5���:zcNv��ߥ$<y�L����Td~�%�AQ�������O���Gv�K�@(:r���+��i����^=�jQ��H�՝�N�8ji��V���9Sy�	`�$���j�?�G��vٙV�p2ؙ��;��]�M�t�4/�y���G��i_N��dhNʓ��g:e���x=dL��*_;���릱k�(P�C�=o)��x�U���-0O*�]���F�_}�x/\AmI	���C)�*��=r��#v+��k���zqy��D�Ms�ؒ�7���'c���
�	p9�� �B�/k�bN!+����8���8��p�:�t�3�v�n�������Ӧ Yr�z�ZB ���/+,A�J%�(P��HV��l��7����6���19ƭ�Q[���}w�[���>�|t	�6�!���z�"����A���S|�]� ��?������@���@O	5�]�٘�^�d���K�b�p�['P�Cp������-h�Q��/����l�����SX�G�~��U_e�vu�7f�jl�㿭�E]���5�ꡲ5���@�S�N���Z�K�N&[3����Sk¸�H�1[�WF�`��F���cO&��:��P�p�[H�2�ϱ]��+�%��u���G���M���Ǖ��z�C���`��2��!��<t�ͮ����{V�1^{LY��
��e4�P%�2����B�{�������߀_g���W���foD��E�},�s>�SL�g6u�Ł:�����W�}�����9h��q��+z/f��C����|MsR�;{\Pc"\�㰮��<�X�`��oQu*5���Q)�)�놠32�/�G������0��<�@
(;����r)�汃>�f��ϮKT򨒥��<��U�Y�x��k��{�`�W?'\D�:��c�].���^��W\�&��hU{�����v�8}��~e5�>�飠�= F��ϻ��3 ɚ�.���C�'��W��fV��)�e��5�R��⦿��g�Y�ދcw����-�he����1�h�˙�@�rb�v8",�P
�A+��|A�4d�oKA��L�XP>��J2�^w!��Af��Ba��F6H`��M:.!���z��H�aA`)􏧠��z�L���Oڡ9�^�h�"$n���(8-�ʮ�:K;Zjd-��ON��:LEl�:Z�HU�޾�>�J4�xyps(`o�o��t�o���ͧ:!S�
�)�%��d��>]�w��� �7�?a7���/|]ӏ�1� #�ߥ�F���A;w�c|Jm�$�X�����{> �-�+A���V�~�w�;���)�t#�Y�_����f���7�:�R��Y5��ύ]�"�r�V�����L+�Q�^3�4G_��e?��jVq	o�J(�J�N� z�=��D*��L!���{\C>S�!�*��KY�6����}���b~PT���3�ӖךpS�l<�]?����r�z�1Az��p)+�
�3�:L��gK ����+S�n!�(�Ǆ!Ÿ��1Hkm"��=��e��ns����߃93
頶a�=���Z넮q*^c����0*���y��i`�n	1p��*��a��iS���.hοS�S�q��o]8�~��.���֐,���54�����7��[���|[&k�oH���H��9Q��;���i����`u�']}[�k�һ���މ%78#�WJ�����dE�D�����8��� �ߠ���W܌��:�n�|��ҫ��vK�`���a�4us�ך�S�h�,�c:���MI��� F=��>o@/�T~��Q��=K�yvJ?!�zF��Ĵ&t��m�Ċ|����i=�FtP��L�	���?�GD~�-���L+i�6�W�\����Ԯѷ�������JȮݡWw,1_�:���v5(�<rF�= ��f�ս����JQ�(X���_�|Ut���a+�����I��3#���xG.�DT���Ɔ��V3pt���C�]�@�dy���ڋZp(��[w�Υ᧥H��V:�r��|6�bǆv9fqmXK��s?��4���Ռ�ƭ�op�4�����Q4Ot���bu*S�3&��F%= !�W����PnzɊ�������+����G���o���1U1����E՞aeԲa��C
Ƈ��A��H&!�k��re��.��ӡ�?m��"/����
�k_
�`0;p^�(� ���?R��\����F�+��o��sG �-�6Km�qP	m�{UiW�#���hmM���55'_����P2)$I=QJ8�&�զ[%���?H9H9�x�{l.A��Ϩ���㩊�����>�']�{ Jq���FRG�e�+�����,��x�e�d�B.'��;�.w�@��3�k�5p� ۾���	F�T�$���9�H�0j���0��f�zAw'ҩ[�<��z"��:>P�i���<˗��&��s�}}y�F5r�
��H�jc3�h��0���@�b0�%x� ���,0A���> C�긢��'��f ��(�wH/�z��_@�WݰJ�@a*� JI�lz����߮M��S�Y�v_Z��YhV�W�'}ͻ{���w{��,g6��}��?���D�%��;��-�i�a��Α���3�:��^�ᶎ�i4�hm���N�rR��Iݢ���g�@�����|bh9���Y�_9��Y�n��
�����*�ԭ�����ZdP�����\J;Pt '�^����*71G�^�D�3�ݮ��a=���,OnX|�X�Z|�e�G�-�~���ܦ� ]�{VS	I��
ԔE��s���f���B��>��3��P^��%	��kLД���x=Ý��v��u�px���}J@ޗ���������C�RPa��Ty��kT��g��iƷ�?a!D�j=)�F�|q�r	8�j����ALa����R�j>X�ֲ����w��"_v�2d�?2>�!��0���~�_�Pz�(ĳ�ߏ����R}vS�b��o��z�,�閠�[4*�D�)J����a��Gh�'>f�P!����_��4���� a끏�"{�#�E����ؾ�ks;�N0��/ؒ�͟�:v�"]k`V#|t��<�KVM�Y�����|4n���0�CԽ[��ۙ���)]B@���^K�k�qK�T1�Ļţ�.f���L�Iۯ&oA�P<E���,�T/5��΃l���v��C�G-�ZN�X��O��\��m�������#<S���Ob��S�QX���.���o���P^�
��>׋G�Y�^MʊEE�2)����*�+�"�Pōt�*��x�O����|���_3Zx�P'q��"���퐢��=�X�<ц�x���%��ezq�Ý�����]��K��e<�Y��d*�j���jbo��ۦ.�2ƽ�0,bG��7^;�H���gA����/�ď��I����Xw����A�7L�j���b�{�H�J��1�x��Z%��L��5)��K97�
ȁYDdW��[}Dÿ��h�$�}���T��� �t�����(�BW�P,�W��]{wyti*a*��cp��D���>�]�!�������!����fTX���mP
�@;R��C�u��,٧���gf#`�%A��"�H�"�^|K���@D��3<J!ɖlSx��|K\�Rr��[O����:8��s���$�Xf&�1Fb2��A�%��:V ��5E}��_>e�O������Os�S(�0+3UY��֭�b�D�Y��CeG.�z���vo��\(R:�m��4ѵ�_:+9���d��TE�~<�ޝl@�*;A:����2��_hr�g�J��vc5�����{ڼT�~u�O^�,�)�P����)�� �>���Nͺޅs���DB' ^��/^��q�*Z�u�_J0���-w��	��Fe�E2�i���5�l�U2��,:�"��tK�|s̠��y��$s�ԻI���b��G�mC�����,�w^?}��ia*��C�����?o�]P���<Z�����m�Y@�- ����1�oXr��6l�S'���]�
c��f�wj�\�����ˇ�V┼/�p���u
p[پ��������Jlfaj�2��e���M�I���\��b���;�����G���!qĶHj���1-�6�	;Z��a�
�n%�}*u�h!��~�3���Hd��6��CLk"1[�@�q�L�'׃��&S�FRAC���h�i}L�E����S��zǷ��� 8��%��b�����U�F��.�h}��S�hfn��0����+�PȌ~I@Sɥ�:<�����č��e�*|�qX�z1���դƉ�6��Xs"VZ��U�����ϙR���r۷�8v��K ��E�|Iz���f" %�f@fyo�`w�)��Ng1�^���	Tb���P��-��6��Q<�C=��x.�~�%�5�9��$9�����;>+)p!.��90��X̝	�0�`�q�Xԕ-�+!df�>l�!�ryi`qֺ캊��&wV)}#k,�N�
�3n�1�]MR�s�s$�  d�.IE/�m�҈T��N�1o&d��LLC"D��[��Y�Br<I!����E��Wq�)]Y�͌��[i˟
@v-�7�"B3�����F���夅�h0��G�K��т���K�Q۴�E^�zp�03\����7�a���y���E��mT�=�h�ZF2��5��EʡK��}$�A�LW*�̲��C#S2^K�\N6 <�t��uT�Y�-W&�N�]�=|�4�&M1��B�f:�h2�N�b�X+c��څeZw�ɸ�B�~��1�C�$���Dp���v��� ֿ�s�懶�F��� ��_��SHFLSB�4�\6suT��u�ŧC�J+eW��M/S�'���������)�����C���aN�:5É=ִN��E�K����䓽�S(݁+���ti����;�᱊C���O��M��]�ܐk ��6+�������:e?�/�	��\d�ٓWnI�A�]쩤�AA��Cq����
���H�p�皀"յ� ��i:��~,�UA�g /j��g�1��$�!y0?&W�C	ѡ�G(	�}���8=U�t?���	�Av��[�~��0��g�OwK��V��+��s(r?#%F����	<LĜC�Ҝ�*�t�;��2�ԝ:��uX�ˑі�o�������#�μf�zŨ��:���kj����/����%��`�\���1�ًM;`\>e
YRd&i����)mBC��T�M��`G��r)�v��?y*�LҐ����J�1Ͽ��*MT�F[(�䱕�vI��w����P���@v�p���#�ᒟnj8���cU�橨�3����'l�w������FC�3(�Q�D�b�7�T�u�!@ʄ�!�D%�<ު��(Y*;�8��CVG�a���+$Mj��9v/�'�{�a.�3.n�?�ǩ^$�M�g�luʧ��>f��P������c+�И������*Y�w`�`�w�WdQz��;Ƀ1ݦ�g$qy�o�M��L�
|�q8��]�P�k����t���������r]0�`�����C�%�i�N�Q*�=Y�"��]	n@8�#�k�I7�5NaN�9|�ܹP
z�๹��<��y���:o�u�/�)&r�-Cr�����Ĵ�Q4T�Ӗ�`�܇zҩ�k���5��U��;���ȭ��o��[=���|��V���>G�r~-Z潻)�e����{���@���
�/��초\����jm~/�A�B�pT͗+����`�f6s�㬵j�~����6�aHH�E���,�e�a ��Q��7b3c�2��7��v+8|e���d��2u�,I�9�F�p"{5�<Uy"bP{�)`@�[<�3���	�Fb��UM�dA�@�b��2_ܒ�s�	b�A5�v��xf�������gݒW� @K������APU�0p����"|�'�h�&�k��И#<^����5!��pp�X�Z�'˝���K�� W"RD��/������q��I��y���@q�C��X�Sҁl��p��PS��oGn�����ֱ�1|��+�I'��7�x���q
֭h��6�kۼ��kK��� I�1�wI�B*wF�����${Gՙ�65��͞����8���Fm�ASk?�0K�dw���ȅ�,aO��F��陀�sl���aa��2HTiKn��ü����	b��O�j���Mo�����K���l�����CR�[���#����+g�ͩa��_J�2*��Ԫ���2�e���i9��[�������%�s8���Jۣ��o&!AI(�:Yv��^���:u�<}S'OjoQ+����K�z@���K�-�	��?"�eU�ap-�<�+M�J��M�d��7±1�Q�P��IAMƯ��w���c+���ơYe5����m��s���<��H���Mrpk��W��i��)<��I5�z�lqY�)���[���0B�O|����F� ��4��5�>
Hi�b�����&<���3Ȗ&�%S���Befj�fi����rU�n+1��y}���H��%���?�-�A����մ��:V��:�<,�E�A��𫲫���_P~!b��y��e����V�(���.q���4
#��"3\~Կ���u�3Wz���|���R�\!��4���;�`|�bՀ ��6�-��:����E�Z_5���y`3l���N-��Q�	�GPG� �g��f��i���7��'��x�}�G3�z|B��f��L������z^x���{e��tV�V>��_�n�)w$�Ёd��y�k�X�{��o=D#+ؑ���{x�u�GDH�H��O}�6�ٴ��:�(o��u�p{G��m{��=��g������Lb�t4�(Nr���$�Hݽ��K�[�E�f���ts�=���m����~�:p"|%��j�T��^Wh�,'FC�|/%�]�ºmhSԕ��u��)��s�8������Ce��>��]�;��t@�Γ������D��Ɉ����<<�T"u	��H���l�$��%��?N|T�m������AP����]�I���bm'�P
_8G���k�Jd�דz|��Ծ?�����>H8~�ﴙ����<T@-�C�|�.2|�e<u��Q,+g�n���Qn/�
#�`0�!�@(�%�^3jO��x�5ڀ��$�3x�:6���,Ѧ?-���xK�L7�Z�Rp��P��������ˈ�m�(�:��B�IF�5C�N�9�bB�7�+e�=����8��LX�e2�=i	e�O�>}��"G#ǉ�����}���:�5�ː�3��q�<͍�-͂8ŷS#�����̋K<$i��^�EL\�ketT�^7�;�e�u��ҫ��XQn����4���8./��.��)�W��G	Mq&"8�#�/el���.*-�ā�z:j���n賟)U�\�{�{X��R�m�*�^j��:p	*�<f�J=��ɏ2�^kz����`�I*��i4��T�A�3��<t�5(���ߎ�T����:�aYaċ&����|5�?�P_U��9_"半#}P��%8/M�pm?�U,)a��/��0#9R[���-�[>gi񱟽�:1�b����z���{z#�ʗ#�+�1R~dp� 0 Y1�O<;1�[��)�}.#Q�ŭ��݆����&�ގ�5���maP���:��k�}b�y�	��6�8�<�~��R��*��+�:���0�� �6(!���B
ujb3a�Şw�-���M}XT�ժ�~��-Mu#���Ò�a"t?u�`
�9=��)���8y����g@��ļz*��5��L3��C�Tn�:wȔd-�g`��l�.�P��c�J�/YB �7�#i�	_�o�8l�+ߪ���#<�y��ru��ݨ7�giI��%�eZ�v��e��/5i�%���GnX����i�Aj�Q��vy���x!B~4���*�?���aI�[Ie;����Fݭ��a��03�Z�r8 �������,�\O7p1����%�!����E��4�)��fۑ��JO���e�m�934�-} ᇯ�Y�Zst
l��4ɏ`HJ�+T�+��H�	c����)�r�SA�,n9rW��a&zi�U�˖�P�t/]\9Tc�WU�9��<�'$��!���}P�W00cq�6��Hl=�f��Q�^;fS����<7�CW7�+9���k�������I�����|A]�Dm/Ռ���Ϊb��lRŎ��و+�"���&<D���\�4�0]Ag�YbowZ�uw���aO��d���}5����݈"]�dz++e�o�Mػ,�!(��H��I��z}@�tn��u���Wg�]�{ YbGEz��})����4t����
#KH�*�BS�G��U�ƛgL!ni�ea�������V�J�tj�n�%2��!{�E2ו&A:`�-d�
^.�O��p�4��UT�"��=f����:eV���2���L;V1 vg��Q����3O��[06s.#uU�@����S���}��S|y���a�vLz�F�H��C�>^R��0����F��<,�C�����IH@e���T��b�<î�T�(��g�)j�[�mw�z�3\ِU'T��8��^[]\�7`�< P�Ǔh�(Q�:�R	�0�Q&Ok�}t{��׵U08�4zZ٣r�4|���	�!dM��ۮ����g��2wxE-��r"��
�}��
Z��'�T����u
n�����V6Μ���1��+��B@��Ba��:Ȥ�V�Y��-��&�^Y����QÃ1ia|�:��k�[��bÛ}��eI��濘y�ʟz�s�����\�%�T�Ow�LzYX�}_}_"���HH�0�q�D;�H��Y������Cwl�;֒J��KE��No�[�N(.��!Y��"�ڽL��J
���L�܉�Z��6Km��$�Hתt��� R��0ӊ��<�"��8���� «w��Q�hr���S�� w���W�K�T�%�s@]���8,����xH����0��~�j�x��]��z�F���.��������dDa�
�9����Vp���DW�<�� ��W|E�S��R6zYF4ą��_�d\�j�@��|�j�}�4��DB�w6\魼���m	wA9@,��l��"�c/�>{]n�ӿ� ���w�PQ���u���Y��Mr��|����;���ŔQ[*W�ʛ8��/̱C�&3�G�U'n��J�֦N�^��IQ=�Y����Ѕ����n�|�R�ߘ̕~N�+� �O��v��g,w���������]uc�g�]�T[o����bCx3"�iY����74J���g�/^i��3�����͛�]����la "���;�(��˳1�%H4�,Ν�Ly���Z��q%�v.m.��u�zT�7�߬�Ɋ���Вi��1��pR�qq����O�s��g*�yS�*c�8���y`,FB���z�E-5Np��R3��������]:��4�$t9����>��a�0ONp�6,�9%;z+�o�7�:�~���S��6L�aOSE�yƈ�g�;����܀'�[�����y�:��PkF�,��Z�h�g@��7�.mCpf\c*�f涾T?�@�6�H&x�����р�[�X���?L7���W U2 ��\y��CBX��ı/����
�E�p��7�af�=�l�Bg��X��������A���y��r'�Q�T�C�bʨ�Z?�����Osk`|���ppWN��1���ː�����4��	�Ι���B�W)�}�x����L- ��d��J���T�$	v�?�aN��r�	��M�R��Ѽ4����湮�Wo�n|�8�l�a��LrJ�� >y� Q�w;��j���:�_�[c�d��[�X��ĬQ5���y_9�X!���=���s&R����u����-c����c;J�js�a�n�w'=�"��	]^������8}�|�L��h�a�k�QJ4�FL���誮5�p���D�����E"Q�*�'����+U���g��Ǵ@|Ά(0� �z!Vuw�]xT!�1��,���CV��ͳ�z#Q����]d��<E����9RH��{�J�}C<��~-�9�ii4�>ũ�n��k��a�����19apK�O&ZG5O�����0c�g��^�� �- ����*����w�X?��Sv�r�Gqdc����:o�)[�l���C��V8�׏����j\��46b���]���bVͪ����B��h����1kO���}A�_#[f��+2 �
��7��x\�M����X��ʒ���e!_�;1O�
�>�J&A�������Z/�?��h�O1	�`����0��h�-Q��V���rFUj�H�2��N*��4@�z��`�~�U�M��sh>#l#�PQ|�*����<��y4�dA���3*�>�f5`w1��3�'��u�̌�v�4�`ґ2aO�a��	bC�e.<+aCi�
y�B,�+�7�0�|wlj3YE��=r�����o�}9��!�^���M��-/T��7 �2�����E�c\#����!����K�Y�i.��8�	L�/���^�FT�:d-8�%�W�F5-^����� ;�c��z���a�7�LIk���Wȴ/�d���r�/��ْ�Ę�
/8�Ei�{�D.����t�1ڞ�U��۟Ϻ��zfH}���x̘�v���v��:t��?��l"�'��N�/�k9�:� K�A\�Ճ�������P�}z�Ry��)�.v g��EI)�DaJ�(n޳��0BH�i�Y�q�63�N�bebqґ�w�F�&��EG�W�Ӗ]��	+Kz�c7��� �\�+�?������a��7'E��_����T�̒1	�^A��P�Z�Pq�)���6�����=��EUF�����۸=�����M[�d9�L!���6��������M��l������ulJN^Au�E�م�y����N�:��<��I���=U��lf�K�����8�f�?��9h��Ĺ�K�7�B���I���E��B�ȯnڗe��Q��H��� �1�c�컥*T�4�D��0__�.RX95�m� ���zu�c���Q�"�kS!*�jO������x)���ȡ�I�a��	G��	�V.��l*r� s�0#��'����\�l�Y��`��K$��N��a93��򹬿�`Pi��@)�#��IX�����Ƨ��d#>�C`':'�Ҹi�E(gw�!�1�+�ys�u�c��(�j���R�g�ؠ�w�B8��{�n���]�~�EB�d=w�@���2�LV sv�2�.�QPx1v�>��z{b����ZM�r)�2T�{u�_#(fR�.o�Q�FR-�*i���0�f���PL&����r�Й�E�{UV��{{V��>S1n6��URc�x�Dņ�ã��T��`c%���`�+��aQ��&���ˌc�X�ASv�䲭�9Z�f·m**n�ˁɌ���Xq�u�l��!zh���@�N^��(�:V�]�}����&;g>��µ�	��ҁ�P'�=U�Tm���f8���FԤvo��+�������o-�"�2���z��Sq�_%j��2�� �,�y�^g)� )��ϪE��~�\�ڱ'ktE�j��0?�ݬ���֙�G�����1_o?���R�wc(��Pw��.Z���O�����*V����Q�p��N
����y�+Wf�~g��E��F9���S��Vz�����6��$٬r��9U�W��3m�ֵ�ݰ���8Aa �+A������z��J�@S<>���z�%����L(�'�h��.��j��g�=��F�ˌ^��n���惦�7�=�V�p�ߺ���We�~%^�Q��=�T��$E��2����/M-3y�D.����_<Nv�y!��-���d�q�(RHq4�
�2H�!Th��㺼lCe�����u}�w��b��q�{67bV�٬U��@�W;@�	-�%�ߟ1�y�T�v��
�����]Ş��|;?�$�A�jT�=aY#W�!����=��!�u��җ*��D�{̸F�[��� �x~@�.�%�c�f�W�H9s�lN�{�M�2��R�ٿ�)c
j����&�C~f6w�
�B�X �Z��]��?m�4��Q��N�H�	:�Ђ��6��!���x���7�X�6��$g<�b{�0H�Crz��~���F����FT�X�b.R�M�#�-#eu4:�]ՀshJV���+xC�J�"���5s ���C��j�Jy  ppX6  ө����e �"1q��#+������)�bo�}�L �^K ��|����p��M�����N��ȒF�t�\��J���*�MܩRY�K1�����C���S�� �"Hy/�����O���>(�
y��r�	d4_k�;H�}Pb�MU��麭�1_V$���$�$v�R��ĕ�ʔMA.��動����0N�I}���n���f��H@\��
Ofy��4���8�"��Y �?$N���2]x���Fvm׻�Im�r�9
Pȫ�T���-�vn���}tF%f�>�0�l_�d�+0��tSL�����3Q'v[��I:�jʕ�ө�:���h=�|�D�=��璣U$�C4m�Fsф�W�����Q.�Qӵ�z��Ov+��W��V�L��}K� t�n��o�x��Oj�ra%���*�G�p��66��B��.��^ �_�6�v[4'�L�I7�'�"��'�	&���o�8DFۂ�{�æ��X�"x_4M��!soM��S詠�~E���C�����~`z��q#.nj���6*ı�qKy���(U%�rU�cW>�۳��ACS�(�'�����X�7��mZj���2�ĳ�J�eLB@DrmhQ�"�c�v3����tF㨲�B�![��Üoz/��5�{Hҗ���R����XuB�%�!x�PЭ��#k�`��.�MO�X�)
�J��и����������x�ِn>l�.�v����l�k#9�Н_ש��[��7�x�\=�0F��6��������~/|j`�	}+�J��ވ��}ĮC�������fޭmu�*�����06h�~�Q�Js|�e��P��H��g����_td�X��3�3��$�&�7�7@��]4�A��{�!݄�:����~�Ҩ�O��xr:�%xMW7��2��Ө����?7[�%�E����d�L�2��** �1�3j����--A�?M{��� 4�_��ԠB��j{i~�$ib�r�ci���Hk°t���&v1�(�����C;9)�"EG֝�7�ty����.*���R$F��ʛ�g/;�����ˀ��Ď�@��In,���"tOC�%����'�f�
ht�:�����?G|ɢS�;e{���v��^z*Ѕ���P�PJY���ѧ|Ȇ	 D���Xa#D�j�q��!����A��"#ɹ��>v���se�����n%s�iE��|NQ��cg���gj�����\��:M�K��3������+~@�0�> �&bX�E�����F�C	�L?a�}�® ����<,��}+���<�B�B��1%1AKV���Ț���Q��<�z�$���Yv��L6�6��[�%��H�(���$��wޝO�I˛�GQ��TGso�� �4ߧ��K�Q���l�2�k�&+��r��i84w�^y(j-���:��/s���:�b�3���Ƨ���MDλ����;��ո
���g~bR̘��L (���j��W�;�����ܵ�J�Md�o�' J�������s��ծ�G�n�m8�G�q�G��D��%��v�m2���/Î�<��d�0�ԷK����W���5uԷ!?H��F�*���F���3�(_�'���EC	!f_��\&9}���1�1ԔvXd�53 ��Z�Ĭ)wҤ�nj��([Q���u c���L��)�tW�LbUȺԏ����#5	��h�q'D�H-���/?���=��+���З�]q(�G����)�o�v(����V���c�,yk��Y�\a��[\й��992�Ƣs!Ʒ��a!���I����G�`'��f��H�v0���������i��O��7`-w�+��91��	q� c��.>��E
�Ű������T��	;��6�@\�p�-71�iK��J@4řQ(���h�*�G�
�i��qJvpT�2	�۲�������Ii�|�� ����sTY��tVc�.x����ɣ�^��$	�¬�^vZwه��[J��a��N�Tk�6��p�p�8OD!-�J��p?Oo�ߟ�l>��*L��^�������&�՜�2�A�Xy4g�)[�	�R@е��co+���Jڠ�z�(9��t�Ḥ���V�&�$���؋��p�\qNmm���d��?������"N��3,C�!�@NM�LK	q����@g}T���M��h�ۧ'��vK�m�n�|�L�� #UV���Z���Ѐ����t���#Q;lHk�g��ê4�ȮS��F��.%w#/�_TAP��X@�l���u�j���^�G\g�t̫�(��Z�������D�(��ݘ\6
E����猔�)IW*��0�����>9�������7ޣ�\����'��9G�QR���݁���hZo�'������;\}�@�#�]�j :�T�����*K~�rt��ϋ���q{�i}�2����B�X;U����̅�U�|�8:��GSFt��[WѨ*�M��2Z^�3�A�(����H�6���Xs�NX�Y.q�46�Z�=��
/]:-�Q'�D���[B�%ܬ^���J	�=��~^.�Ps�b��9��5�Wh7t�f5��,ޞ���?�����e��5��˓�S�J̥;ۿ�Gb[�@���_}���dF��p�Ŕ�̑�Ց��*���f���p}!��/�\f�ȶ��n-][��ߕW�@�r:5��I4�xO��Q��Q3>R��S�x'���Mۭ6�5,�	p�8]�Ӥ���F=�`/�(S Z��ӥc3[���FD�+U|�����w��B��+^������W)��o˗*� �}��������4������w>�㟜4����w�&a��t0g$���$/A��[O�)�ƛ�t��-D64�\荚�'�d��VNx TV$���^z&[6�`�U�m]�.���[�716W�z6��C��-�A����b��d`�˰�� �Z���P߭��m���M�6�%%�<�K�l�7
w�S�k����IP�J���/Nw�p&ϫ�r��J\��ƍ'�����բF��c�e��)W0v�!�O��9@��ɕǵ�Bi�K�t�{]��|�"�ӓF��KC���l{������v�c��K�3�g��$ή��0��l���uN"�C0��So	?̦u���G��*�U;Ƭɡ�B��gg��R��(��*�zv?���"\*��7�߆?lo؅�$���hR��z%��TO�=I�^T�1�A��2n^�.-�|��=� �zd����p'�Փ7�Ab��(���O��"�!N��ͺ�tZ���K+�y������'zm�}&��@�`C���t�v�<�HP�\����_Ԉ�֙�T����eN�)EE#i��_��7��K��\�NpV��)��C�q,a�1�Б�(6,���l�2�gGxWo����(f�\\ wsK�W�r5w��^v�D~�4,2]���>����B�r*�'n���cj�����y?z�����W�y��ksaq��+
���M.�ZdSĒ�鉃i/���]��P��b���Z6zz�}*�hqa|���7�|C��-���񗂹�� �)G<�Gw�)���ʰ�nх�Ι��Jq>_��'l�Z;�=F��5R����߀���ֈ1�v�扂	N�1�aX�D�L�:J��<�8G����z
�&NU��V�ˤ@��=�0��4*<Q!��E�/x'�t��-���uB�R)�ͻ��E��]��g�؝�_�4��@���Kk`�����"����fUȻ.�@��M K��O�����FQ���C����j!F#z������O��cT�	eD���Hc�Zc���"M�CJ064�-9�ק��m�~�y��";�5�na�s��.o�bR��>P��A���̀>~��������Rĵ�*2����V�`7��<F�v|�r	_h��=�W;1��[2&5�B�0�?I�F&6<j�Y�9!�Ƶ=�	B�2�U3�3�8�c��"U�B��	���U��h��[ao��P�t��ؗe�p�N~��f(��^�Uu�.ALt�? �R�=�?��u�,��A��G����y�] ��[���2'w�$@TR��+��3O	ڶ<!��k�G���s,�f�|��/��(n���_j�����#�v��8��v��c�d��P��_Q�u,�������狺ww�bxƫ�ca�l�D��a�+l�ԝ�f��m�B�_��	y��_KIӒ���ވ�S��%��ʓ��bsZC�#�!څ���Y���y�`ɿ.�������'�
���כ�@��w�v�T�*~F5�l�j4B=��%.Hγu}j\�f�h6/���M/ V=dg�Cq���pdey��4ˈ�"Z��Y�ա��9�*��^}f�ο#l5�՟�<{|L�]=�Z,_��l�i��n([�����>R� �U/f:T���KQ���-*��򺼨G�;�0�sG.�D�x���I.��V4t�g�e�-3��լ�zg���@���Gsou��pw�)�0�Í�{��>󏽏�I��D��Y�S�\t��;-�����֐�]�n���2�+ye�f%c���żu(�D�tY�]��\�aOɳ��'�i�|y:UW�؅����#P?�Mq?���f�}ieY�gq���ICHC���v��M�P�z�|0�_P����s�nz3��E�y��g��wGā��mV����t���l�܏��m���a~�P�t)��wK�]�w�uf]���TD��� Έ�d}׃���\�v�Í���E��uq<��CZy�����9 ����;��RV�Е��3'15���"_�B/$����;��> �*x ۠�W/��Op�A�=g�7��g����'���� �^;�ê˛�`��I��0�'����{V�Y"V/\���n��~꨸)a#!B|ܩ�bmܬeU�?:���	�uګ��n������dP��u ֠?˯�HÛyS�� W�J�&�P��ݗ�S���/�,�_�5byr���rJ�E�/�^O{��~LIC�����h��p���'���ir��h����@�s��g�:������'~��|V�S��b�pa��ϗ#+#���C��v+1q�S0P��C�}5B����6�)�=��i��q��8���6̍x�@�G`I	�_�K�#��p��8
�9�������?'�
�X� �O�?TD����T)��f^�&p�f��$83�+ݰ怋�Q;�|ُ�q\���ܸ�������/�Ձ\�z�����wםf��e���m�;ql���,���]!^�����y�,�G,�oy��jT6:���W|��X6�ɪ����]O�O.��Y�%c���^�H���N�c#��]�K�Bp����2�}N{'e��b����	����&A����;�E3nb}�s�<�gU�y'�G/�T�����$���eo�}-_쌒�tY\q���(7�MdҫL��_��W�K��z#��~X+,�rk��sU7�T��)��A3-�mEv˲p�Ť"�Z��z������ݭ���GJ�p��:�x|>�������^d��SJlV�]�f��MJ$m`���1,}������qQ#GN.��&���B�(���8B�8]�����u����.�J~@Y�Wg��%�d�5�͹/\g�$��T�h���=�9z��}\�!ͼ�~����#ث^,��!�0�Ҫ����9�~��A'#u�K�"e�>�u[��S���ޛ��xdݠ�ܒAdmB]p�|*#w��C��3Ȩ��T��#��/kP����Oj���C���55��`���m�	��nA�J���t����u|(z�$;�&����}~#�����B�xZۣ ���qk��_4��o����Y�ϵ�В7^�Y�y�-��=6P9������`�'s��Co$��/Qs��Q{�׶ ��������&Z�p�D�	tR��At6�uNJF�誈�G+�>ΖJ���wW���_�S0���6�_�6ly��-�Q���H�������Q��`�e���^��J{$���8&���8Z�e�9��l���S��&Z��Ki1n�����Zq�%�=Q̢뼆E�$+�3���A{L& n�ގ�,d���G�8ܲҪ0K�δ�aX͕��~m��ְO�r��^�Xo��M܊	#�R���s��IiHGv��h��I��ǬiE��x�͂�ŝ/��Vz�yd�a;x[�.�IcR����XP4:������|w���k�`�Ooc�ӆ�}�
�N�/،����	���f�C;���"�	ۃ�{E��D����wћ����@�=ٷz��4��g�
�Q�\k5��G�<��o��lJ�!�p.�У�9�ӣ>;dO1�$|'�Sy|�t,�.*?d���L�WX�*�� ����o�;.w�F3bض���"X�ߑV�k��p�$h�*�0T��3�D��#Vk*��6�3Kv02�m!�����d�,�]n�x�� �y�8�.�������]�$��_���}����0�<K���{�����v��Cڶ�%y#�u��QQoT<��@Զ��ON�0�UO��b�^|�b�s��tܗԑ������ϧ�&�}���:]w�� ���uV��]s`ScT{��7Ώd�a���F-e���ia>$�֐;VN(٤ �Nq���9���ύx4U�"H�4v�%q�&�`�=]��FJ�Tu��]%�vDD℄��ޣ}rQ�y�mև*MIv���쬙��h��t��2Sţ���i�M"�_�/��S˻PH���"V�2�^�\^�uH,x3c� ��	�����*
��x6@>X/�I�M���ʢW%��)-/IH��{���ІP��$ ,]�-{d�H�!��c�ש{��¿��d��������\:���q��-سf趁��c�,`	�y�6�6g9/�}��|���-�cd	z3�St�K,j��]f9��VH1E���	W�dH/�����!��|�Μ�^Ֆ�'Xԣ��[������F�q*i������c��$�]���,��$qU#ȿ��f/���,X���s�k�7]��)},Ҥ�x�ɥ97b.��V�g䮷+ :��~+ijP�\�_��WD��l�G�ˤE��";���g�����WB?@�����/�0�MV���<Ű	c��I�Ho}:A٠����@H'�����k؁�X��)��<��@ �4h�����93����fo��ow�;���`�G�O��Y¥N��\Io���4-=*�+�"�@F��*w��f���5�
�a����~���T�ccƊ�m��?�������>����F�DA�}��]Z���BN�����KF?�|�!�1��M��J�d6�}	�^�6AL��g��~	������P�� ������y�Ïf�� %��������OV���m��	xN��� ���/ tʇQ_��`��R�Z�ܰw�=��T���K�|����4���q�����E��K0'�	k��ޖJ�n�wf��!Wx����4E[�c���w��O�]H��Йt�L>��0���B�>ǟߘ��0�}�b�p����O�L��M��1��&Xj�*k�U�F&��DB2E���%���^(��6�����6q�ޱiY֊�8����OJ̥�K�QM��K�$s�~mu�1P$4j�#����GѴ�t')��>�U��ۋ�����s�6y���}Q6'cOz߈L\7>X���S8A�����Q�{B�db�T(�h��j�F�;�d��|;��fTٕLρ�����
"��>P�,bj=}�e����C~�e��H,���W��M̧��KI'��f�:��,\�[s�qP-�FQJ��'
��������;M�]�>!j�٘�sttc��}+#�{�[\h���Y�1��:�cd�@��Yԭ��ؼ�+��~��׾ � {�~�s�S �]�(/ruh���h9��ъ��ң��8��p��̤�p(!��[Bj�*��*��l~�*t��5�~�	Zz����
/��E����b���(R�H�k���^����ղ��0�9JI6��l������9O�-����Q.9~'	�C�-3p����}iࡊ4���F5)F�@�vߥ�ni4����F�����=��o���ș�����q�^a%0S%����1�f��Gx�C�S�-�]\ȹC1ԮP�8$I���O�DY��
����4<�^5k�+��UV�@�&h����B�����;�N��n~E����N�m�tV��a�TGA�;~$���q>O]	�`]��x똳䳫���\aEV�y�򱔃�tn���J�+��g�r��eO(�����j�G7Z�����O�z����_b�����[�8�A���ɧ����yL����߿MĦ��Kb�^��mPD,���}s�x�������9@L�g#o/���!�S�l��G�R���M�!����G[#���p�[�cQ�QP�b9�s{�p�^��3����K���gS��(Lͩ��0 -��ԗj��5BR�7Nd��⁑
[�)Ir�Ջ��@c�tR$&���{�-�v���S{�D�ك
�X��zLp�ل������~鴇��/#E���̢0����wsc�������b�a�H��ғc~����oȁ�~�z�Ń�,�|�$�)FVB�G�f>)�T8�˭-P�@��v��f=�f.�X:�c�r�
��pl��@�M&�,g�&�>x���Ք%וN|�2��)�zG������i	��N�
�������B���1��nP�A��Ƈ�P`��8�^=�~;*2���l��We9�����]�U�2<����@�b~�Z>�|r�{�;�a���r���ٶu��,!H�Y6�)��v뱬}�B
[� ��G�2���8Q~D,^�Q�I��d�\�ˊm#�+�|3U���ל�Cw�,%��o����5���A%�;�o-�Q)��������\N>6�x�}�X�_s�$��P��nөq��0���	)�?�zZ��O>�E�@ٱ�[��x4��WiP�^����M���n���%���'�A	B��AΠ C\�7���@�r���/\ ��v��V����� ?��W�O��d��'`��^A@5��,��L��d����y��9�����4?/�+r[sK�B
�8 �+�ьL��2J$��l�8��ֳ�E�-�ok�]�����*�0ў_h��.G3�=���jK�k�l��Cq�eQξ�S�`+��d֨�pE�4�����C��"�:6�0��~oe���⼨͐��9q:��y�l^Pѵ�|I�۽;�X����P�MWAa-��>�`��b�B%'솔��')Y��l�gZ���9 ����唊�T��J�;K�8����ծ��L���P�����1'�?)v{�W䃺�-..�h�u�U1��z��9��PY�'U>{/�:�	A�������l��<C���B*�n�ɡy��c�x�7k6	?��h�Ș�6=�͡���%�j�Ō�&CEۜn���Xc �.�"��K���@�zQ	-	h�U���sWf��b#*���,�.*��9~6��Hh���f���c�SO���Ȩ�u�]��`��_��ӭ�@�~���_}��Җ.�(WmfS�H����x�iKh���ep���龺'f���p2������se ��a�"��8��'��y����/��H�LF5/-�� )�.7��	\F6�~���������k�v�ALX��^-�-�X�^.�,�9
rRk��j�ߓ$�n��5&���
�S�4��]?�vr̭YL�,:�r��-a�k�rW,7F"M���Y��$l�@��I	�)7B�[?$���r'h=�54_��i~H�1p�v9��2�g93����(
�ӫ{���*q͏m�'����CA1�!�ZJ����>�]�����Y��:��>9l�WY�x�bۦ���kæ���P���$0�/T�<�(DvB�B�u��_92�`D�4[1����#��)+hZ\��u��<�<��F����"C{5��������������S s�u6�����+�7��#¬$p�.����(}��[�`⛚��k��r���+R��__��o
�\����/0 øڲY'��+XKx��S�p�bxc;-%E��6�~v�9g�������y�����x/(��Q���R���6���]ܕ�����@}B�|@�j�ٱƋ�C��1�G�tR ɇy{$�j�m�k6�JG�7f��}���6X�	9�9
<��z楉h��G$s�ݻv��(���V���U4%� �(�&zt�m���g��`	)[���=��3�~S^�n��6�u����/�Hw�ޕ���u��i�A��׎<:�-���hb�y��:��:/�23�'��������@�Xd�_�
��;-��a>��h� �B�q;��M�qT�*l��b)�婙t�XYG��ppW��#O��=����u_q�
aN���Z
�§�&��qq����!-ԥ&n₺J��~���e,�AUϓi�]�ߵo�NYF2^�5���*�y�MX�Z5�X�̎�_�2��_��?��.��G=L�6٬{L>�J�eo	�*gA�k�����{�N�V%C��\!T/kٵڰZ���d�H�r�d�-���Z*���ڭb־)�[�辎�������$�>
b�K`@sG�:H���"A�$�<�֌1��Ӭ�Za���(H	#�L���cN�*L$���$)uL	ֽ9*9]��fs _^�������R~}AO6�"���ST1��{�4�P���ں�p���%�R��BB�԰2ʾͻ������s7���B
g�H����L���_�>�x�n�6���y��2%ABr�yS$+�)�].�I�y�A�u�N7�?�s�M�TM�TVVʊzR����f�6 /����*��^K�L�;u��-~�V�d�u�����y�˧�������R�>��mB�~�|�>;1��c���$ ��+kv�T6L5��V\�˸e�季�5A� ��'�C��$�*+o9�z������g�n4NH͇�խK��	����E�Y���q�عōA���9�Դ��#z�����Ԅ�]�Y�SCzM�`B��Ck�GY��X����M���f��n �fI�K�a� H\�M�K�xq'5�u,Z������c�n��r�Tlt!`�v���9Ox �;#�0ip�V�w���a�o���<�|�A��~�*,0G���`����F;�[_"T�h��M�uX�4��Dh2?Hzƙ�у�I��D왥�[�;��9Q�E"Q�j7~mO� ��{^�����G��.o�7|���6��-i?���@�fm;��)�Z�y(칳�3/��ܰ�m�����AV�u�q�|��e����Q�h�!KT�C�DW	���"w1OhK�_h�������!a#%���h�gˈ�	0Y���'4]�lL���3]3닟'��v׃l�iV���R��)�3���)���6O�2@����ϲh:T�5�ئm>�2������&?�|�F� ��p�-���h�a��a4'Y��K���I��0�W��IM�L��K̀�Q��L$����#��e$��y��cX29��ۆ�[7��]
l.uh�P���zo�|�����\o�Q5GU(���/��|c?�0��1^	7�?���r�3�	��ŗ��ⶩmo�yĹ]�Y�s���$�g@�)5ޚ6޹���4��4ԝ$�g⦵K�DLż1�v��'!��;�b7���B15��e
x��Z�ґV>�IԞ��I�=!6Y�R/k�z�b�� ��&#D�av=3�yٝ�t�o���(���4��&�@B��\���wl ?�u,�x�R���zg萡��{��)n��xIK߂v�.����Sq�������~V�^�mE@�[�E�3N
6F�T�I.V���ć$_.��n���[1~���ic�x�4.�{�-�X���0�IUԻ�����]_K��rMS�KUq!���?��+6�$���e?�" ��0	v��273w����c%�T�ȉ(f;f�ݪ�w�M"	>���CO���=�qs�f\pc��(���`֗]r�F��E��3]r<<�A��R*^:[<-D���1�m]diuFY K'HCvТ�AG��쿺�]w!�D��-��񲽹��(��8���7�|�v�J5��H�3��M@t��ن��w
�����f޳]�am@$��\�Ŷ�!+�����Ѕk<"嗾ߋ�bm�S{�1�
���RE�B��U��VƖX�\����o�ٽ,��/���ı̵�?���nr
���2�/ǐ4aờp��f�Dt��!� �����j�i�J	Ǔ4~�*��~�88�״�I{dFȩ��C���	V�q�"J���`�'e�j�
M� ��Jc0�=�p�}���i	���̆휔-aVā� �.�w�:?��|9�#J�w��.��DS�?PYE�ɤ��i3Im`�z��0����1���f6O3�FAr�%_� ���M���D�"��Y�j��b�����M��r��̺7�1�I	�'AZ����-��'����-w��)h�M�2�.`>���K�|ȝ0�]��#���LSF��E	Ƙk��(��t�����X���&+�dL����f"\5c���O->�g�ї�<2���䢤hť�̢�<�L򹼃�R����n�V�}�������+�4+:��x$��5��//�oQv�#�F�bȻ�E��G�:>6�/SW�t�*S����n�/rQ��"D$���v|��~.���ũ3UH�j�t�?�y���)S��,̓�cU���*'���M^U�f^)�O��F��S7U���\�m%�Z����*��4mm�;
1��JK�]r<03���3�lp*c���=��H�k�S�����ާM_i2��/&��< �[�o�����ʖ�v,��76�H������o�3Z�3��s?;�%u$�6�mȱ�A���j��!�]J9�]�#\��K�X�?} Ue�JL�+��4�/OY����"D��VE��撅��}c<=�?ښd�4G�|�A�\�n�A�ܓL�;�U�?�B��@P������L�����p�~hN}��2�	���⩣f�������!`P�{W̸��V�I\�!y��X�Y|��e$%;��/��)���^��T���������J��@��]7G#�!��|��pf�b��I3Xt�/(\��G�}p��r��a�W@v���p}��_Qm�t��٫������~+�:��#�Si��4��MW�.
�e#��\2%sJH�D�E�o�y��\ӌYߚP�������K;�r1�j���i��t�{{�Vü���q����葎��%������p=����u�oÝ+�9pGCvl��9����Ws�����Z�Z�\<!'��2L�8�,2���u�݌�7��kkNRYx+V����<���,1��+��8��u���_Zj��2�#�q�t�څ|C�rҤ��@�';��U/bT$�y�0],��;�YE��>�/.��ܸ�A�G�d��5cA�{-_��݅����(:ҥ��b�V|UH��� �>�7�4��z�&�!b�TƸ��n����w��Iβz��J�Sp��FI��e�+.`�Ŭݧ-��BA��Wl�a֟��!JãJv��٧���Ux������s푀���!u_��nHw4�޶��M�JH��J��Խ��X�i�}���P�`�'�Qhk�Ô����p�a���i���"�Z���8U�W��c+ϕnp6�8������j^��R���r�;�D/7�H~�S&ţ_��c�'m]k0�F]�=��J�C�3U�E))o:4�1ɲ�wi��ʮN�$��%�@[�8ְ��Hl�M��~�Bփn�e4���.�F_��*�&Ef�T��LR�|�����;/�F�zZV]�i�a3M�AH��|�1pKLk�RK��; ��}�O��E�-��i��L6al����ut�l��^�T�K��F`�gb�U�ؽ�$ǯG-_�w�;^�����.`<	���d_)5��8� ��Ԗ��>CkWYw
�	�t�����O`Y��x��@�AE8��L�8��u��r��,^��ý��.>�礜��k0�
l�0�vj��(nĤ�,4���Q��]��Ћof;튓Օq��赪߷�.ǥ��7�82�+T
J��*���x�[M�+�pC�iå��E��k�F�����#~@�0!b^���a/wZ�t/Pp¦c�V�| u��o:��LnR7o?��+͔~�#�*0��T�������s���-ޅ�R�AE�=��ΐʹ��,��yT'��kK8ä��ܸ+�0?�q�4��$?��{5,�%��M�Awk�~�{�#���.>Q%Gt��&������|�G��IK$g�nP�c��V�"��\�ua�U���Bu��\�9<���M��ުG��!8/ [d2#}?��5|'�؟�C)i:7����j��A@�X4�ܪc�1IG�y;��_*\��n�:��욝������-�c?�ٶ�c�����^�����O������U�K�TT�r$�_ٝ �3�l��pX��N"`̦^�m�����c���,�7��-�!��}[��i������k�I�F��U����z�k&~�/���_:�<ȍ�m�%��G@�jYvL���ٗ�<o/�՝������'��Ԡ0��s�V�	<$Tӈ=ukf�`i���:a3c/���<x�(����0�-dMV�𽃐�Oj����_~�[t\B*ު%o��j�v�񓚷(�g�h�o5���;"�)�֚��u���ݗ��	����F��y�nAh?�c��rs��|l�<�c�s	�ܤ�U�~�3�K����Ž3?�7���*]�>�%�$[���܆���������*�M�i��/�I�sC�T����Zf߿A�Y�����ҿ��#��{F��^��	\�]���SD\qU�'����֜@$�e�(�Q9~�ħ�G��˷V��+��2^S��i�fÞS��|X��!�}���9(N�ł�O����N�>D%v����8	��PJ��v]�Ll����cH�Cբ�:r5�?{:�A}�8��%�U�K�$��R��9���&��=���v�ܪ����N0$�XÞB�u� Ot8�_�3�-zp��]vE&�4�*$?z�ٓR�i,.��`m�B�E1 Y=�>��R�Wh4y1�O0��`��"�j_}�!� ��e�����YORr����}]���a|ɼ�Q��.�X1z���I��hXC�ʻҟC�|���X�0���M���'��^�|^�}[�	A06Z��-d�'�N���hwwy��'ҰƤq���1T���@�)L��y#�	��J��M�d�5f��N�g�F q�u�1�'f��۫�sNΝ]�2���>��%��>� ��+����'�D��/�X�e��1����1���z �EQ~_3i�x2�8�UF@����bB�ψ˰��h��0�|����%蹙x�t��7�0p��&��_�>�qW�Nc�IA 1�Q7�d�e��.��ۿZo2�����Q�K+;	l�D	<^����~}��y�����9���(��4��݊��[=���9Om�P��	������E���C�r��=x�c���dM�����$EU�_V}"��a�2����߉��n�ٙ�.�)�$#��F�ar3@�m��d]�'�-�V�ϟF����M]�۠iϵB��G����}��֍��x�ı���
K%d��P�f�zDY�+8쐙b���f�6�e]�����Y��F���k��]ɒLZ6�5�Iǽ٩ �>��E���˹�}h\=�dwX����h��%�s�6�>��u�ʒ]S�FX�K�;n;���Q�`	$A�43��OC5�w�=�>��⳻�S��%׶ l���p�ÿ1 �'cK�$�q��#��&!\̊^k-˦����M*-�4Ҽg? j�PDp:m���7l����b=Y��W�
�Gl�o/46%y��Ǫ����2���&�t��J�t;��- ���݌0Fn1��y���6�j��e��i=�(�ɹ��JV������)�wqt�J�<�����/a�y.3�V�����%}���!41֒YZџ�@�2���9(4�l�ΓT$���s����l
�+V���$���P��e�J(���C�WB @��駊�D9
���A
�vZ�Z=�XG��_�*��m�(����`�&w xeo+�T�fm_?��f#�y���_-=���4rq�:�(���Ȋ�0������%�j���~s��(��<x��_1<}��w�{��Q�_f�6�D�s�����)i0��;���)&�����3i:�r�-ePj��aY�C���ٯitq�WlѮ����pW��{
����Si�*I���.�Gm)��/�5W�Ymq���)u�s.�p)�2ط{���Z1vfzX����j�'#.��!=�?0��i�XY��L3<h�q��.e�tj?��mg@A^h���b���y�-����2��Z�9�\����X�~�f=���x�Uб<�U_|����j�����Y���[�߲���o�"�#�a���n� ��w�~�
����������x5��X�b~�(�������⎇L���A���jTKGv����
�U�����L'/r9"�Ȳ��G!Wu��{ʝ8�wnc�&�fnMf�۲G[2O�<R֤���ך�篹{J�d95�x�H��1%�+�A��'t�;�{��֋Ond�`�o
��)}]���K����UEI��E]��8��"`�hB�#��������hlh��@�[iaH��}�};���:I�gZK��r�O�o�oKׄ�{�F&���~?��9�w�H�Z��'�5��+XC���":�&g��D�z*3=�9q�R�H�̀�?�G�ſ:��0�k��uƎ��@�Z&��MnͲi��h(��፺������s�}��.eMAl����/Ɓ����t��Ԣ������$ψ�߹x ����DpN?���UB�ӡdzp�B��^XnR5.�9�X�%�ꐸ���,����u�xހʓJ��� ڮ�	7�Vt?"G�0&�F$s3��C<iF�J��e��X��}�	`Y ��.�Y�`�Q�󲛹cz�3=��^U]}�Ժ��#�K@�!���yw�\�
��m�}���0hK�yȱ�S��wm0�q�)PsL+��캀�j�(B�R�+�4�#�I��¾����j�]��ںh�J.3�`K��Mс��wL�Ӏ�"^�}"���YL��T�p��VԚO�K��ࣞ�x�r��+��-�l�׬����Cf�"�����c���v��f@BR���;�������r�Y�n��l|6�[�(,�k�Ok�5e�mh�:�iӁ�R�,&�r%�9�y&�yd�s,|N�?B��$�NY�����:ᬝ�!�K֙��p��-R ��@{�����G��
772r��bvyf:5��ty����"IH4�*|�刦����5�[��vo��\�n��~���lR���<�C�c�6�J���k!r&���u����:�	k)�5^��U�@ŷ2[��',��BP��-�1��23"<������z���#I?��7��M˛��y��Âb�q�$3����_�w�_酛��	39j���C���I��f_^'��yƿ�:���ҙ;ӛ��]��K�mfe�q3Î���U=6�f:�@�l��^�~\�����u��ɦ�I_���|��̑�pѶ��J�YL�L�&n�!1�v��Mg�\D&ò�S���r9VT�g�|/�����.��3����3��T��Oh�G��K�#�+�ۑC�ϧV��[�p���/�`���	�S����CZ��)��x�	2�@W0p��f4C?�`J�� IѨ8þ	���M� Ͼ��
�S5�)v x'���́�����e ��V��!0���\��$4����u5���	�7��23j�.�p��8���8L���e��u��0���@a޻��Fx_��<qH�K����=Hÿ���5�l.lO��V��ti۬�	�}�A��P�9���_�օ§�e٘9,Y=�<�%^m����j��d�&n<I�aI��;�rܨ\ݳ��O�u�{���U7[[z���E�i(輙��V$�8M��2"���Eӊ�"/o7���7���4���Me��d�bBP�7������zg��Wρ̐�oI\�֎Z��/�4�I�Q���~�Et�@h$46}��/]�d0�u�\�l��ݨ���)>�E:kE(��.U���S�c�����S����C�8�$�-h��i}"�����xil��"��iܝ9]���kHJɯ�ŝp���3!Ѻk�p}��%�����,������6�iV񇪞�!���x`q�l ӻ�G����$_�5�l��5���]pS�_a�ȞlFdQ�8?�g!u��,��	��h��(~y�"� �4몚ŖrH9�24?hc�L�ŁDa�P"kS�?����K��=C��넲ϽS,ا�����n+�y"ZOPI��A
6Wb��Ż��0���������W����K�������9�k�����ĺ��C��iv�����j�Ml�F�<N��r�������-'�R�!�l�&juIX ���W6�L��, ]*^��L�l�l����2/Eq*х~��k�K�J�q� $#R<+(D���ϣ �N�X�0ڰ�_�,��B.�8"X�`7�� �b�@==�Co�D��_�+���e�b������2��$�%�#%΢oh(X#{#R�&iG���/j�u�\z/�=Ƨ����5/��H���)	{S��W��>^���a��v`h���%��)׾����Qz��[��	��k���pz|�֣�d�O� 	7��>���������u�����������%�%V�Y#ޕ���|(/9B\��{|%����R";
i`��veJ1�X��ȳ`�@KIr�i�1s`����Y�S��H�)���L� yJ���1m�z��ml�nAS��t�յ���3]�V����zgp�9�a[%�r3FN�wҔ��XߐHL3��q.O��/�c���z��bWkI]���B�ék�V�E�Έ�]t��A�����٫��
�B�p��)ޅ-����?�1�I�l֥����zd�RA�0���݂�(���x��R��p�@�d�2�G��inh�~��u�EL'y���G0�`Z��Y_��C��x��WP����S�w���k~��aN� ٺ��$࣫r��0&�/樽�nB�
�U�V�^>Y���}@ՑR3��s?�~�(?}�(���{�{��>���KB�D(bQ�1-;���#�)9��m^�4ΰ��K�=A��a���_�]w�q��ڟ���G�y�*U>8�pS��:�I�O��[P8XVI�*��x���9u~�S�?��l�A��O~Eu�T�i�8�=�G�G�����1���lт��<��$#3��[�m�^^����o<�=L����FX��X��-&4���Iͥ&��Hղ�3�SsV���6B�C<<�	�L֯��)
ͤ�U����2�Ci��e5\�XJ��]����"�;����ｅw���I3Z����05�"� [va���k,��.qW��$� �ݾ�-�2� ���_�]�x�7xx��N�z�a���8B-A&Ib�	��X͈����^.����qKK��t1ΰ̇#�IL=��^%9����mq��yr�ﭳ�ys�.-	!���6�d�'\2��A�	f��1����\i�9 9c�i�&d��G���4=�m�3� =�@�����@��W�T��t�c}�r�dX��V��D~�y>#Eg�l�b�8~�+�
������qΈ	~�$��'�@��؄W�1�:a�e��N���3vSb��,��L�@��Խ�z��r9���N�c�t�� 3;!ea&�%�u���-��$�as�]� ���K'��_���1;�-0�0����[��%����ox(#��2�	ONlXt��4�|͞E���̀���K� ���0�:�tX�#��I����iY���c �S�Km�kAdHu�E����1�~����rh��	wr�"j��:}Ǒ�2#��Q��Ł�M��e]'�� ?d{���Rț�q*������Wh[�!� z	m�J��\�?f!� WEP~)��k@�f�g#�}01$U�Q��VQ�_����7G,w�l�,3�WTu��9t����6�{H�
i_���6�A�����"�;��e��L
VJÌS���gM�t�Ր��^�NQ�3�X8LM�E�#V���EŚ��2đ[�V�xh悈�a��H��/�J��X`�"鼸Y�'���9��V|&�7������E
������l11����Zg��M��p<�y��G7�Q��^�<~��V�n�B�ۗF���)�f���U�h��`#����>n�|?����p�E@��z��q�6ǜrr{Nj�.�F�~4�����`��ɪ��C|t���-0�Q_@�#�'�d2͕@;H�1�0V�Y��k��bi|���F{��Y5�x0@�%��>^D9���;,*��r�oq�2�l�5�Mj��)��B�?�^��Bpc]1Ի�6��	Uܙ��?�1�b��x&��NOHv�3G:�g��:��a��v���h	�q�H�È��Q��@��+Y�\�Y��� CM�I�G����4�:]/^����A�3$�H�߰`�+��Țm��N�4�U`1���/��c�`&0mT�=�hڇdI���,�d\����	�����ttL(;+��S,��
@�i�B����b����$�Π"���mjz�3��n�W�p�A�|Rc68�Uy��賠�>ե�iԔ=�z�����݈�q�X#��AQ�W.���!A��V?)X!���� ��D���Ȩ�6��cb�����I("���)?`,�y���\�Q��s�����m+kl�6O�G�OA9�/�c���09|q�]_[{���m7T!�f�}O3(1X#=2U��9��K`[���L�U��N�ڦ44d�;�9b�{F�e�V+�!�ê*�AS��D��AAP����(M�PI���?>�G��yj�����w.n�E���8/����� T��g�B������X��c��2K��S��3d������q}"�����z���r}ʐqA!���t�@a����Y�]FLK��b�Ip�7����O�)HΌƕ|F�*3-�J@ ������7�~���bZ�?$��2|iЦ�.���8��c0SS]^��m���B���e�ȇ'�_3(e_�՘���g�"���D�u��|N�[[�������-��Gq꼮Ц��'���Fi�z���hK��%0	o��{4"1"���r��7���$8�dhK�w�5��$���kD+ø�����|�^�*���ٽ�@ZF룼Zxt�w����q4���sgR��]�.���#����$�Vd�������B{���%���k8ZN�(-A�qh����>8����5/���k���}��)�-9��9���V
�U2d7�z�K�J�[c"�٦�������PT��
�J���,��[�,��E��6���~�U ��?W�����~�>����0��%d+<��>gN�R��Sb/������M5{1O��Ԁ��Z�+L���Q�i��C׻����lu�0.O���n����H �D&}Z�^��V�#�gvٳ���`�n�{�"c�������ۀ��S
#i^>l��x�#���xD"��1�\�f	s1\�g���KO��n*QE�t
�Z� ,���EU�G;��mm�Sx/C>�W����I2�/�h\�%Ҙ�{�C��f!'S6���)���VXn�Ɂi����Lr��<߬�Im��S�����T�:�%<�AȬ���T󻡭�a��F�&�X[�p�PW�뱌BgC�*��oBi!X��1[�-�sN�LrqS�Un�F@�m����@��W�!9��N0���R�n��;�˱�a\����kyэ���)��H1���G ���T阥:����2E?�8��Tw�z�T0�w���"��z��
�GA������|	T�v#�!�[�z���s���%�A4H3V�JG![���ZJ���ɧh�ʝ���Yn��NsM���x������Bd�X�������sOg	T��Bݛ���Um,-�u�S<7e���X7�����٬���8� �����X�A�+�'���+�nl�a��.F4�4����$��)=�!���{�B�4�抁P+��Md�A,� ј�J�T�x���ʆr�e���sf�۴��ǳ�i�@by��ALo擡K�Bv�5��9%�K,��s#&����W��@�Ts.�_�KS�{���'�I5�ħ�9��(J�&�<��c�V|�@m�.�OֵjѝvD������$-][1����>�:μbM��1�Za&���1���o�e�;��������E��o��o�"��o����a���Y)��B0�-?B���x���ԸF8���RX�xh��1���]F��j��r�X[vI��Wж�ƶ�ܳ@)��ܵ/�Vz������ ;ȐN������A����S��Z�g��5Ő|\Q�<��p�K �F�V��8xߺ�a��ex$''SRH���7��|�������N�~[�
�	�J��+0Q���>/+u*�]W��ظ�(j�~y�J�+BX���h>I��q�����(�碾_��m1-Zm�	�G0>=�P�����ѾL��/��P�P����Y1 ��5�ϱ��>r;��zZ�ϟh�4£�����Qq�T����)�kR�����^�����⡛��$m-�/g��0�,�jT��?p%]r�Q�tG�R4���-�X��hnG�摻t
/��k�V�����n�X nP��w���fbj,n�j�R�P��:��%)��q��� )f��G�iA@��z}���R�h��~��j�#�H� ���eO߬U��N�ҭ��|��#>b �;d~)�vH
1ՄK1`�÷V,İ'�N ��ǭv��NQ�m��k սD��+�y������:*q<�e��ڽ�R}5�$�!{�;,o居,�� �yW��93Z��rk���DK�x��߂[��.����>��νqP�����B��d?e�^�T|���8]��?�*�O@;��0�+���%ϭ�SW�c&f�*��C�Di�� R�+F�0.".b����i�J��#f0�9ul�a��4�
�bҪ�ֲ�jJ�A��!�ߋ�C�hi�2�O��q�q�+���Ӧ?�lU\SR�<JW=yEH��=����R�#�Dr��Е����Sáwv�+�8��c/��7�md'��'���"�Tf��B���D�Y~��Vָ'�&T�=:�۝���.��y���g�Y����2.�'&={̱�(X��`�g�3��)/��Ԩ g9P��w����Ѽe<����i��۩p�A��dO{�vp>��E ��e��"NQ�XA�N����-�WhV��I��=�h�)!f�
��ABc4[�M��4�԰Ow�"�ܴ۟�l�Nr��T0S���0(Z�'N���_���s�� 5}@���?	�j�=$ݼA�n�H��/�k����t����nl��XI����D$���mb��r0���q�fy�"�a�|��8%ޒ4U�'�F���t������>�Qh A�^�Hg0��{k�w����u�N(�o��~��E�G*g���O�j�]8�V�̝+J߸K\��ǫA�j�Pif��Ni��"�_i>�s���t�6
�؂JV9ʻ�Պ�b��`4�������sX���W[]�DQ����\��颅�gz�bE�
fCId<Lwi�˖4S�Mm ����B+��&��/�����ǒ�2� � 
5���Z��c�����y�P�3�Q�]��{ �uv�����S�Ы�n���ye�6�LeO��I@:2���l#@���e��2?�G�i��7m-u_١�^�6�s�U�&����<1�S��<i6Z᤽iT�4��+	�2Eg�Q=%�?�����=�~�E#i���0(�չ�j��KO���W��(�0݊#䈘T�8jC�����e���Ӫ�x�(�!�p���)_Pˊ�+��A��&4�&���ǎ3}"�uo�c߂�n�>�E����z-췪�����3�y��7JD����5�f�\� �F� �u�*h5���3�2h�J������@w3�Z�D���p����� �:���F�Ic�t�a�P�a�;�vW%���zj��T�Q\�K��
ajK�?��z�^��ͻ"D�1n��_�hAuj�v6��uB�yw�����Z�}����k�u�]]�_�k�>9��tp\[Ǘ��y�s�BAX��.k�7�b%C?d�c�/�g���g�el�YV^'J���������an���@�;D���%$IN����k��kw�t�9�F���,̔j"Y�k'w8���* �֌��������qsb�$��޼nd�����,,�Ȅ�ϩ�/X� �&���"��~
-�J��B
��=�#�r�ӗ4�ı�+���>&s�k_=����L���������L�C,�'.H�-%��ݟ�#����i��w��I���g��R�J��]�(��t(����8�hf�l�d��u��o� .�&��{g��T�����8i)��H�J�12�~}�<����ׂ��>�n^i�����W���A�R�M�Rx�rE`EU�U���ِ��޹e,h�3R`��K�@��u/<ʲ�š� �ұlE�n�˪��X>za��E.Zuf$��YK7�������b/���`��T�?��у���������n��|_%x�����x� ��Ւ�nha���(ؿ~�C���	��� 9U��>���߿�l�9�'��WPAm��%Aw�; ���+v���|1�K�iP=~D!4' ��]���Q�,�k�ƅ��=G|�����k�o	���"a[P��Z<��q�a����G9 L�zw#��7J��6����ҷ��1�/X$����'5hY_��E_VM����|�����u�k|c"*�Z�D)"�͟s����?oK���J�Wp��Pۦ+O�l�H���[�6q�� �cd�&�����ww��;�~��F���ߺ(*C�e6^p(��t�����IP��s�y�d��"���)8
���za	�R��x�t�*%�5�t|� ӏ�0Vs*%](��ma�?�%daSY{���gh��0PI�+m}����Ӕ|r��9.ۼ��;wڪze�2(!�.͢;3'#�с~o�󍉼bH�#��L>���Q$��A���Ҥ�r]qq��R
���;ZA�
�(�'\R��߱x�cp�sd�ɐm���i僐�#`Q��5�s�R@�����s��V�$�cŝ���l�ԙ�=ܳ&\�z0�p��V��M~q�o)-�u�����X�#�.��!�Z�"��y;���Xj�C/b-s����Vf�v���R��lLSƩ��^�D�o)㋣c�/�y>S�#Y��4G�AU9WS�ls`���y1�Bi��}����?�D��l��L�p����蝗&�-�a4q�y;Ε�q��2�/3A4`��^��^���ȹ�I0jBP���A~���=<2��
��;Q����G;B+2i`oZx�S���0�
�|rW8�c�^�*�����^�ܖ�@"��d��o%|�p�����X"�>Bpl�a��Q�Q�)|[X/z ���x��O��ar�`��I��&}.hWNiy��{98��p��j�#�����X$�4���s`��Ea�.I��F�Q�M��p��ᄩw��Gǈ���JO{��IZ=|�{�I�q� �����3I�����]�Έ.����,�ط?�M{.3.킖-�T�tF�XB���Rk�
�	�%5����w����puߧ���/޻a���6[4���&��O'�lp���v8��&Q%Ʋ�"1��������=���Y��xce���x��W4���z?���8��e���.ֲ?��uT�]P(�v�=�d��G�W�f�iF��iYP��%py�r)�Nۿ��5iFS�.��$�$������mnz��[���~�vœK��YX�xp��J+�w�=6�&" �\lh�����:�Ů�����5a�����&��v^P\X�-Oݜbn���v�</Lf�!�h�7O�P�#V�>z�H���fD?H�U��3qŔJ������y��&�Y����oI�o,��F���Fj實�%f0L�_!�s����d��%sM��IK�1���I.s8ꗃ�|��+��r�7��@�S�w�m#-�G����7�35�.��X$%�^�cl�=����s��%"@>;�l+$�-���tt�X-�j�m�V�.����;�z��^<�I�	�P�o�g_���p _��d�o�%֧z��!k�	��r���xG0O�k¸t��5?�a��9���PtI��7���;�`FQ�W1�܇"�u�f9E�zGl��!�N,s�>�\�)�q�r�K��]؈�ّ�n<�/`�ޙ��ʝ>��`럼n*B��X|&�U�&j��m��u�˲��P�|S������]a�h����{���CJ�i��#�4�]��y����U��M	P����$�S�m^jM��Ҏ!�î��� m�y~�v���uԴu�
�"�,����~ު���	�����D^t]�D`�K ��z�_�Q�.A�x.ޣ�{R�%߯]�m�Rj�&�8I��[+3;��-��h��r���YA��m��f�����~�^�_9��s�K�`2�k�B�Gpmq<���[���э�ԗaU	�°������a�jF8�SJ�޼�	XW��t+=�����@�M%��0JH]�V�.�bzlC�f%�^��<2.��k_�d�-"�vQM�LNeZ�E~f*dTg	�鉮K�!^e�?UJ|`C�����"	s#]^�5�p��h�:1]Z̬����B�6��G阻
͏�K`��s\2w.<��V���^F�R�cD/o(�*��O;>�1�S�{%���ȧ��>������3�D8�J�^�|M�������M��������E��_�CV�o'��"�ٜ�{.� ���m�6�E�.�靊��OW�З<y��ibaV�����+�}���+or�'�� 6��J,pd_l@A{1�2:����1^PzGS +���\|�i�#�!T=��b�c��sC�l�a��(�a��d2�H�+�����l��@���° ��M
�mf��,���������8O�������0=���1q	5^�k���߷�r	�i�Ɨ��x��R+4�:��L��]&V��<(ʉ��Nn�ɛ���i���y��(�Ύn�~ �`�����w����3�,��ơ�[@�
��U0�G������о5���
�����,�.�hƦc�[��,�-�6���F:��BQZ��CS����_uK�]�m4�3�c�>���R���S����W1Nc�*L�|tYׄREui��4�_[d\�:(���䦓�yB��h! 4g���߷��?�����O�V�Z�QC�(�3?�c�`����K���m�" dd���FϨ]+v�K�h=���e�a!�Ø-_����1fQ��\My����S$8��6k}��0�|%��S9k�l��7BP�9Z���؃�N٢W�ؽW�H;���5U����,c"k��aL�K��%��	a|��i�'�Q\6ŕY���FkI���; �����(W�P<��44�7O���CC]˩�r��Z�&�cO�6	T+����-�Io^p�K�\�k�i�pc2��X�p�cHk��ڭ������j�79�Lb2� ���e�-ߏ���Z=�o}D��0��1��U�nړ��?���M"�^>���8k�Ə&��Mn�k{��Z�S�g}�������!%u���q7{#�8��Z8긐=6hp�B�Q�1�n(����������qk��8?s��H!"����~�w0�,�X�0�zh+�t
�/����am,���C����䇋�D"��/���m:�h´��pS���
�QKL}���ViZ�c�H�q	�q'���]����/�P�?tF����1j��͈�� .�yvF�j��a��!�1>���n��o6#�1O���-�����'��^�!��Q��Y�>p%&g�:���9r��l�q��D;������1����"֝�L@g5������d����o� 	���Q�t�!��Ď���y���V�J�Y˃6��5���X�/�y����7�ǖ�v��n3��ݥ$%�ܳ���c���Nn�m�V z4�x���ɾ��f}�h���U�+���*�Ё
`�t��a-#Z~���ײ!7�&*��O�Y8����w	�{��4����+aua��
��#^���/�ɟ;�f�K[�� ��*��Uf�?Bm�&�-M[�,�[�V+L葸=��k�+���,�A2������D�&��hͮ��.�U��4I�e�����co���Ɉ�����a�PH�Wc̏ 9�	���w볌kR �	�5v=��+>�A2����7Ce��t	<��۳FaE�mp*I��Ԕ-��տK����m��ZG��� �~����(4�sԛ.*GG���n�&��O4JJ<��_�f�d���+�c��b�J� ��7w�����e�/���L1���4�3��-̸	=���'&��	p��4�Lw�E��Y2�t��Mk~v�K-�؇K-'����U�Г���C�M������Tµ�Ѹ�$��=E��t���� ��}6�%Pn�m��C|ry
���O�����t��~\"��LH]}s8e��n5����Fa7�LU^˷���L61H���UV2�&��&�I�m�e1��1�<&>F�8O>]��s�8얎��8����i(5~/^��]%n�j"�`�c�#��������]J_v��"O1��eZ��'w&"?�K}$t ݝ�I�uءQ�[�u�P%�ٱ�.��Ji�$Wc@�4�3��%�����:��Z2�Ѷ��J5-f$�T%[��M8�G��������̰�	��S57�z�iF	�?��f�0����h���f?|J��?狡����	*�##�����{O����$��U�^e�}b2��Im��r?��>���<���ӑF��T�<��p{tg����,�9����9�R��(\wY��2�`q�����uh��ᬑ?���{��NPg=)Vȃ����F�������:��)���×�إ�ϔ
�{��w7I���l��@~s!ڮ^)�,d1���A���]1����|+.0$�����Z�IB�/��?��Voc�NRld��U��V'0������R���S��~�5�C�m!���>�1�<���r�F­�+�6ru-��??�ڻ]�_��$�#ˇoRa�E���Ńړ��)2L���}��o1Q����wY��t�B�SE@��K�uF9I����,�y�.A���^o�~��B�ŞPU��kW%,�&׎�7>�g��M�[s�]���籾}��� ��
j�v!�R�$� g�x{��~�� >�K(e��ŏ3z90W�Eb��d4��:��[�m���'��q�%�Ĺ�N_�X�O�Ԣ�RV�� ذ%������=��`�����"�߼�Fŭ�vey2��\u:L-�"��<�:�`!l0Ԍ��{������Uf3����Ϊ�
�0��!�.7*Kɧ+��#_�,2�I�<h9q<=�8]t�M��7�9�t���6|�������3S��M[Rr�TJ����*Q[
�g���f��g�VFa ��}��h��L�*! ���8�����m�F�S����|T"G�],ށ3{[�������i���.)-�1��PǊ�m��w?�xN<m.&�d�Nwq�ڞ{À���M����Y���-貑��<���Yϻ�==m�d���KF��p/��k��9�KxwUmv��W���' ��_�� g�dX��I|���4"���8Y�"O(-C>��~
B7 � ��e4�H�kJ�>�֟B5�w+�}�4���Xܯ����(�RƮ��"sj���O��TK:�78�
�?*�k��R��6a�o����t��ڔ1]��}A
���$�3�^�4j	�K��:��m
B�� y�a�x��A���s-U��G.�;��,�^1�<�P�{Y�(
x�?9��Ӣ�4�*ꕀ��]Cf�8(�:�_�@��f��Z�虈��%���z�� ����rذ5��8wX=4F�y�)��DD(g[����@sP��z��K�E}����6R��Q���."�3T# +�L����B�)a[�r&�4�
S�I�&_�l�֠�{��uKulm��03'�Y��Ѓwd��Z/KK�����u�R��^#�{�(Lԟ>��%�ϛ��7e�c�1�K�.-�9rهFI��0u�����9+����~u��:x�X^�L��V풚����*�Ѧ����)f���Z�۲)�������n�:uW�R(�MgsĹ��'����j�\T0V�H�؈�&ϊ#��a������C�9H��҂h��z�t��R��Y�!�;��
'�e=]��i�6�{����X$��F"6�j7K�	H���p=�S����}��:�_�Fe�[g�K�o0�Ngսg(� ����r�4Ω^�����\[�^~7���'!�n����\�)d
VG�ڦ��e3�΁��fх�����Ф�%��QI��4�&)B�6Wa~kkHE��k.D�g5��.d�Q�^L)�O�}U���s��}�n
��������F���i������/`ƴ����ʉ�� �pc,�\�pR�r�?5���;nwI���PD&��ʦL��o����|���.BN����������ɋ��i��d��i�
R�n��{ |\D���)r���O])	�#��!��T�Q��^���ѣuԕ������r���N��D�Ď���b=��t~����KM<Vi��cc�i�d��>�c�u�S�(�`[5��U�rx��u,e���_5�<0���B8&֬�:�w����wnQ��N�kf�f!*j�I�)J@ս��B�qK���-��5�������m���<*�e���#���)���n��3ȻtS��JΖ,�c���P��ytƓ?YsBga���@}���}BD�#����	��ᘛb����I������
t�%���5�������E#����D��VV+}���3J�+5s.���w�w�H]�<
��E��!�V�Wu�9j�Y��-ա*(���W$QckT�����Yx%t��	�/��0����aWݖ�f�����!�<�f����P�NM}���Z7��<x�j]�Y��i���o�o�o�TQ�2��n�*6������s+�����9M�u\�o�+N�+`\�4���O�2��ڕ�By��7q���#�oD���d��Įܦ��5���,�.��h��RA<�MC+�ll����d��	�dR�<n���0��Q�%O�cB������652Qd�q$��j�)��f���a�Pq&<V~(��rnwDP�2˦���_�hY�o�#��$�?�)��א��=u�QZe$:�w�y�ӯ�B���	���n�G\
�v�����̷�v�Dwt�������1�)���S7�")�t�*�}5$�6�"r�]y�mg2�<��i<%3�g���8G��CB+�Q ��H#(#���<Z7��#���^���s�ٿ�6n�g� ���O�p��o3�m�ᐃv(c�ՏR!��o =�{Y�CTnְ��?Q�a�1��h��όZ�	�v�u�n>�3��\�6��Q�K���ӆ�8��Ǣݠ�i�~�K�����#Rnkq�[5S��G�գ]EW�u��䖠�HE����Έ��$����l8I�;9��oN��{�#��qp`�^���'(�v��D����F�"�']�j�1�NT�<��O&�'�|�gӍ߈{�]��.'��v.{�I���6��^�4�#j˖�eGѢ�����W�����@Y�=�l���jm��,5�t���#��e�^���'f�+��i�ہ��gY!��M`�:�$*Ǡ�7R�	`.+O>�W�ӑ���ח@���C����M�|�QC}�n��.U
���h��I�2ީ�W1�E\����"�8d�_a��rO9��0˵݆����Hh*�s�.��/�^%�Z��S���$+fH�@q��nᅶ������ү����ɠn.i��b^�9c^��+�Y*���/����7�+V{��߲#�_C����rM���&Nt��^�u���^9e}����G�g��?�
��L]��'\g�
�B�G�GV%���>����I����m�f�g��w��[�r�)@(�F%�:%��E����
%}sv,ż3��J�� ����E)�$S����bs%�7� �\ʳM�v�>_T�|�\�{��7��t�-�m�5�Yu��p�~���`��;�J����4%��F�Z��""K<��I���b�zP�q��-��*p�8�7닇V��p0?xl��g�\�E����a��\���\�z���?:F�޷&r��Y�%����~r
PB>L�(�ï�󨌫�>��N3[�LT	�ɫK%��.�uW���Q`)v�k5���U�?��x1v�'�	<�N�R��tZ��&B�3u�v����F��<��|҆�v=���jVEWEC"�� f�.�2 �e{���,2��`8��%\+�Ȝ6�4uf�z�!8W W^}q�R�aY�Sv����_�7 �l_�������WX5W��?��m�uc�+�)^^��z��/�Vo�����Ȣ���x$�!�Q&���	El�sF[��L����SI��KF�jo>!�7�����>.y� ��E��pt&=Ԏ��H��5En�Y3�"i�;���x�`��S�:��) �ZJW{��i'��B��TC�%̋0Q�n��{�Hꚗ�f)TO_��:�h���3�1��֔��Z2�Lg2���|��[��N�a��Xxz��c2�sA݁st@�4zk���\��;tH+4m�Z+{�{W4MT��(�?�h����l�?0qg�F	���FR�oD��GH�{:y�q��+sV�b�����I�N<�aJ[�{�B�mj1,�.S<L�,֑YV��y�J����p���J:_D[T`G���&�.�����1r��&��DC8��:4��"Y�T$XD?����#b�f����j4��J�����)�.t�����7ځ��^'y�W��x/���q c��O��W<˾{i���Xu�lw����<#��&s��$�D2�ì�B%�����1@�U�G+���&�Ǯ���ٮfA�Se	OM1�VP�2�7����;�Ѡ�v�=�l*��R q�jNMI�=�Q�[. X�RP�J�<�����t��p�	�45�A�$Ԝ�x����p�|Uk������\�mo�6�ڪ��"�����L�ŷO��0���&��7ry\�����Y=����cg�٫G�{w�7�<�9Mvף_�4_0ygV�wV�ܡڶ�����5u:Fc%'a�ˏg�H%_�2/b������ʔ�ѣ۾[u�1�q67�op��D�m�#d}������Q8\�����Y������^���8*�t�̸@�C=)M����,V�����(3�?eS!9<�Tju�RW��������*�k���1ڪ���N�$��_�*B�a,�:�m`��Z>��س��'k@s1 ��U}�R��]�C����(8|��g�$��H4��D�A��n�i�k�e�4�[���:��e@K����iiW����)d/�cv��yd����}@�������E�I �m�N>�
늌Id �\´�_[��y�ȫ��T�\$��Qe��,L�/��'�ICa*�l�5�6�����5"@a��B��V4���ϲ��N[��R(>�#jv����IE=*�Z ��%���櫖Ny%8������˒r-�Q3�ļ�)�Khfu�����)so;�`���ў�YӰ��+j��M��GcD�V��>��|*@<3X��J@��0-Qp����V�p�J�<�I+̋�ѓx��"N"����Cm�����.��du��4�$�`A��6���
HS�2�0��Ӵ* p}��vI�������jH�I!4s[l�^ICX��1Ԩ�^�hk\�I�r�6���S%p�� S!�����F#lr����>��ܿ���s,8�Xs��[3��s{�<�c�A�Ù�Hˮ1ѵ'�g���zi�_��599��l/I	�+`h���4�A�;޷�P����,zA5��3If�1/`�FiŒ
�+vq�c���F@�l3TO`d �ed^�.����V�"}c(�π�M�4^}��[�z�%�9���j+��i�����S�mn���Hه.�X�xy�^�8��a���v��l�ԣtzX)�]-�A2��ᤰ�N_���j�%��9�rƈs���KH��������h>�E�>�W
M3��So 48dU��� !�P17���e������+o�ir�"ªKKz��D���-�LS�_���`L�G�U;=? �^�J\ԝ����o#i��]����( �t��R�"�g^Zάm�ҝ�x!J����<wS�-HU&�����)�W/b̷@�_�O�&��x��2�/��n�$Q)��N����j�>����}�iοh���N��#�Hp�n
��|�)]?�Wp��l�y�ʌ�C`ݤ�~�A��%���[���бy��� ��x�{K��`>x�p�Z����L��D�ې��n�feE��R-%���ւSR�9��/�D��b�ae� �����4Qta��N��R��Z-/L7���E���t�DTQ:EN�t�XOU���A(��r��b�8�/kOV���X��!ت��4uō��k�%wa���%�?��,��;2�E=Vx���<}� {m���6|ŴN�F�A9��: �A�@�)}���a��U��%m��{)o�dr��ą1HJi�T�*�=Zy��Jhqs��jYh����`&%�ܜ�[��*%D����I���������谛?��!��|~$�toĽ��]r��5H��GfI&G�'t��%� �2:���J���5�M�_ ���`����6F�}1Q[C�X��s9��ʴ�����5��e��^�L��ҭ�]'~ 2�i ����4�݋�VEv���̘�z�4�G�1;]��<��p���A���!:�6��dyv*���DtΕ�ԧN�p�W6�8���Y������W��k�ň���Ia�R!y0��%�΢��
�_�Uej/ ��Y�qR֑��Ũ�W���x�bEز��aɞ`�*ȣ���YZ6Ӵw���Tݿ�|e��,VF��^v�r�_ؔo�A�������&y�����]���&� �L��EɕN�)��A�@Y�9�t� l�6�]\rf���It�<�ZD��U�����o��H�l��������,b����K ������G�+����F=�59A�"�,��%z]�5n�zk�9e�a���C0vc �1/��
 `׽h?�Q�Z�*���	c}1JJ�%�e-C_�ph!��7�e��;�|F���[泌t�N׈:��%k��S����aٝ4zp�*?��r1�0�+8�/�T} 
���Y:ϭ�d�$����ͼ�m_[�"�j �[����t,S��
�2���yNE(����,q#�V�-J^L�� $�{��
܁�$�B��~>.1��^#S���B�A��v�h@ZM��>ܦ�
P����){�^�ne�7�{r�ÎYX��,rX��<�1y��k�Y�+�|����@��;k��/,v/�H�����X�����}���.��A\A-�i٨�&����Z�Y/T
.�甽$ ���!�����ʆ�=��kSy��[L��ڑ�g?/	�s�~�r����BNDA����ۊx���J�����X����k��������u�V�j��C���8R:xs�+RЙ2e��`����Sg��D��$�*c�&o�N�qڴ�6Ԭ*$_��h��.����w����|!p~�s<}������Ù=3��.�|ah�,a���7>����>gS�:�/D�1���5$���
�5���i(�]��u-�Ԅ�=�!ǉ��}6�)�>`K�j�ƏX��uB0$�4~Ԯ�,�?)M���K�#��!��oe9ku��'Ik����Z29Z�z�l��&4az�]z�v�{xҐ���A��]��@��4�v=Nq[2��%3]�e�`�&gF\b�R���>��{&~><�Z����T�w�^f�W1���=���0�+GF#�A"!����ؼ�&���*�Y����$���\�Y�3�ĺV2;�� )��Ӈ��#�W2��iCH6٪�����֋��z�L��*S�H��d�h3�sg��!(օ?�x�8�["[��s�}u��L��<p���o�������V|sye]Zx�{f.)x�=ɪ�+`�&�F d��3C| ��1i^����]�d�&��h�������̉sߠ�� ��Z�]��9+�}�N�'g�K�g3 )"�mz���D�4����0*�~:�������L몾������?4��LEA�spD����ŘE�VEU�G�AMA�4$���y���?���9���Y��}�v~ri/4M���L�`�:NL�BE�<��k����k�Gl�3�z`��	  ��&��C��(���=���u�$h@�_�?��pYX�2��eTC�hX�Is�넕M_S������Ɉ�:�c�-�pu��C˖r�B����j����U�j3�����d#�0de� 	�`c�#,#��S�>�J�hA�Щ)�M�g,��F2�j�1�d��L�Uz�[���T,`�w�����Y˂��)2&/{���n�t��Ԧ�T1�\ɞceA�p�Y�P(H�eA����P��Ht^�R<���7��]L~ѡz�t:7x���ڇ$�=xׂ��[0h���������Q��f;K�:�\v��Uؠ�7H�Ӌ��}�|!q�yj���H�
X�9u(��ח���bĪ����Z�K��31���k���8-���U��rv�7�$��Y:�5g�".£zX��F0���i���JlRx�Q1,����B�M�2�'wab���P��_�.C�|sm�QL��ӝ��D���%�xԜ�s�gOȎ��ս'��� *�l06��B����8O�t�������R�z8�aݾ�MdX�^˛�	Qخ�:'�E쾕g?���-�dϞ;��_]���`P��(=E 筙��noб%�LEi��f"˕)��8#��;��n�B�"1����Y��,��9�~��S6�+1����P���� ���Ek��������0�S��e0�H��2�.��V^�y�
ɠˋ��!��Z� ?��.8���A����!*�ِ@<�1�I�v�g�׼�Q�v�����)��p��:ʩ!�~a��ȴ(�ܯ&���oȰ��F�����Vw�b`���j�W����c�!Qٽ>�����^W�0�
�p)�R���h%���*�r"�eQB5�� )��x�b��R�a�dkwھ��/�l��/Bn�;A�ĵMgK"�_�H��q	|D%3���}rF0�r���*����J�hI$i�d�A�W��i%&J���:r^4؆��d����hI���ҨN�='�Ɖ��)b�'�K�J�������I͛%QZ�<gp=C�����k��Q��%���e�s���#�����I�<�-�����}s�^��:�.�[���3�O��hf1Y�n����oA���/N�P��U�x�s��f���ֱaf��{8f��TYT`"p��`bt���ÿ;N=>�8���YwT�<�c_���d�Z����E.�I��f�/PѶ�BuHt�m�����r)�Vq�|�YJz1���������|yC���	� ;}g����]GiC��#�f6��p?�ڽ�SWhq>�4�Kp�}d��l�����S����0e�2^x�?gZ��z�o��<2lP�M�h>�dKa�.�MarH�ʚ�`�nPF�'/k���Jp�e�!K�N��{')�[J���\�猙��9d��K�L�.c�0G��[N4�a�J~��̹|]AD�UB�����/nqCcf����Y Ӎ�ÎZ��E���O-�^E�tW�Af/�D����ᓁ_�No�'�q2+��Twy�g�I����U�}M1(
rPDaB$�iGĐ'?�qs?���|����6�p��� rY4b�ɠ�f��>R���ͅ���P�	��$���>�5�H�,?S�1���M����e��H�Cio�tP8$�2���ڀ�ˀ�ЭŨ%��<��a4�@{��/8}��|[��%�ݝ���!_m��g0��9�z�l����򫩌f#��։��俼%!�;�}�9�5�8ⶢ��k�6�UC9P.�J;I�T�ɤ�Ǖ�{J>�W�����J>!�E��ь9����I�ѻ|r���z�هQ2��
Y?8y���׊������j��ujB�ޘ��?AklvK's�H�&�k�2��N��̔Fk��5	o�`$�}>�b����	��/�u��x`��d�i1���}1�F>���2N������*�o�y��3���i�X��Q�j�/�~� Vu�l*�>=q�YZ
��ա�d;_ұ��.�wC�#aܿ]��U&�0v��u��#y\�?�,"(��7{�,����[��6p��e=+tOF��y�V�'�6�z�g��6D���u\��� �~�6�0�p����-P��-%�2!��:$Mz���!�F�&-b݈I�B�
�_����<�Q|���U=���)p�Ǵe~xjl�N��2������_3���7q�zd�'����
�ˊ��u�D	(�S���^U�8�>�a�"���K��TZ��I�(-s|]���{\�W��>d&�)��XJ'��X6�[e�'�y#�O��z:���������E�捌����I�$�	�-���)U��y��� _j#������ϒwVv����&�f��
��= >��p�����G !��j�$��5���jƝ�����]��#�-7�gC3`g�M���ǻ��$��`�}�N�J�ϩ�O���VF�����&�PD� oV��gn0jf
 �d/���+Pk��	�%O_+�e55���(����0Z]�3�ڳ�Z	�b
���0��Oߍ���A��!�
�����!�E3�H<�RS�u�*uK��s�\�\�5�ixs�A��H��'g���,�M�U^C��������`�+����~���L����/��h´�/�~M���/�f�A�p����~�@� v8��B�M��/��X�+�}!�݄�.���\�^p�D�K�γ��c�2:îS��x(0=N�T�ܙ/�U�h�����K����n��v�d�� �Q����\r���B:���]�q�i����E��+�A;��]�Ha�T�ب�[m�j�C*�5� 7P�{���L��W����"���ILj�wy�>u�k�z&]��b s~i���u��u������a{���Z
GસQ���W�r��N�o�Pu���/j\Y�X�HF�3��Ma��!M���lN��CL/��C�a���j8$�kV�?�}�Ђ�	�Bd�c��4yg`���h{�5@[%�綝�~��ٚ����S����zwy3�{�)��Rr�4������/�Za��P9�	LHZ/���	�L�M�P����s����������d��X�&�r���O��Y�aNe���X՘��Z�0�U�Cg��t�c�J�PҾ)]����Da������GO�Iuz��3��j����x�;g�,��!��,��Y�"e����f2�V�l+�P��[w�h�'-�m�IO!�(K�Q�����N:���fR��@��R�"�lǗT��x�#�f%��t�����4̠��1>0w�q�Gt;R�lDV����rDo�+#J���@�*ڞI��D���AD ��D�Uf\U��|����.O%�Hz$�@E3��2�#�Gu�-�ef�To.=��M��~O�K��7<�B8Z��2������C4��
Ⲍ0� ��l�>�4ö_�
Uvh0Y�����G��^Ĥ�T�ؕ��o���3T��>G��L��ղ$���\��G�l�>X���B��W��8y�N.������G9��E��1X��_B�^N`�ƛ�x��GԄ�$�U�k�y=�; - ���0nuc���I������}j�$�Lxi8�J��1ѳ\\baՖ�������
yY")��F�ր	�PH�3���˹i�l��j7	�	R��W�Iz���=��0��z雵թ����.e<�����L���-�2׈�th�������z��g
���;ֽ��&;��T#9�9W'r? d������0)xNg1�A�:)��l� ����∷�H6˿}���܎�YuS���
�3�M�k�i��"��a�ɿd.���2{�#��s ˸b05��}z50����N���t K�d�:Bc�. ���Bww����}�[�5g�*$;�w�������v��C�Eu�zp�XUQ\]F�\��ŀ�M|�\��e�Y��7O��f��!rR�b8��ף��"�X薃7�b��9���baƆ������Ռ�A<!�.�7��7���QxR�[TmV��K���fq;����:���=���r�k�}��Y�<���CՌ��eϱ'� ��fp��Aϊ���G�t�
��/1�5*�~Կ|�pڐ�wo�J�#��L)Q���44����ǡ< FΎ��h{��%���r�����& ��:"�aC^�m ggU��;�`guTn٠��sJ �mᅙLM03�$ܙ���#�b�E~�95��5��Y�Q���]����������B���$NFH�<�S�u0�<�M�ܵ�{1��A]6W�af����[��j�N�~�<H�0�
��;w���+D4DX"�W,��~&���S�N�Y��3��r"/V!��Xw���y0B�WH��N�~J̷ ?�� ��\�.�I�L�bA��!Ơ�����t:<�`����p���b�j���{��>Pr���,��⩷��pЭnq \&ʋ�-����J�)�L툆��ğǳ G��v23e�P���^����`�x���d1����*�9"����n?ƕ����-W��,CN:�g/G�\�:��M`"\�(��t&��DK`����1���_S<
�p���z�r�Y`��8㲶��N��~�h�)�W�+E��]|����x]��iY������Z��S�
��~����Ԭq�1�./)��xm%�W����j�&ʱM��Ui@�fK2+��y�]xYE��FaC�z�����n�-��i6+Z
����Rj�EΞ���2��ػ5��R�v���7���Jy9�X�=m�Π�ոcƿ�� �������Ek�5UL�7-�T��zh�J�.a^��r�Y�����@�fߑP�j��� #�Pt?��g�#���B�^����|�{a}l�]���?��U�pm��kB̳U��3�J��K3�����k�-��-�f���C�ٓu���Ih�#�]IQU�I�{ 7��:�p�d�z�3b<�>��/��d/E0E�c�h~TQ�	����r?7�/��<��8�k
�gN�����t�������vz�D'?���A���NO\��-U�{A�o_]}�si��S�?��47uɡOVX�1S� ���6�j-��w܃�72��gk�3��>L�mg�r�� ��A�� ��o��EI"�R��>���
�:.�=���Bgo�|>S�
�3�|(�Y_Kt���dr�B-�ѯ��$���\���|����D�9i�E����L�^Q�$n|#��M4�
[G�1dا��Ʈ�y�>_���l8��5�^�����wm��>hߑM/�!�%�?TF��_���2*���%���

��g<&?��i6�%G�i���Ez��=��Z�Xj�ʤ�Q�y�^d�V2�?6����ɿ�k�&q� y'U�8K�ݾ��J�r�q{~:l'���֯�k��8  ���'�C"P��M���'JpD�`�x�u��^Dh��L5���U�����q�9%����$�&��c��|��L7�����ٳWc��Pv	ߠ�)�ioK�Y(Ml`��ȅ�5�y��������$D�V
��v����C�['�T*7`�{��R�|{��'��ƈ�͜-]�p�99�Ht���)�����k
{\��� ��߯��ơ�H��g�ꋉ؟�wD70���\2�ڷ�(�>-��+n=J��e+u}���	9��z|X�sT9�.����ͣ3���n����f �㕀�4�C?H?�[q�5�ɠk���#����񩘯�A���W�����ᡞ�1ǈ�$%z��p(M�!���蘏�~��Y�\�5(�x�õ��;��I�ӂB�m��Y��z����o2!����۵���M�����Hl`����i	eA� Sy܀�]6�m��gM6x�#�5��~k�
�r� �8��6��}"Ttq�",R �qxL��՜�
�xgC@-�44�F��H6��QZ�7{&Fb�֭1آ�U]���q��>�b�ʋub��FtKT�"C"F>�eU��|,^'�����ًB9�>tei�mbt��(Wt�Z^�]�堸����1��ζ$m���f�d����vD�>�y������@��|����2�w㞇T-hqG�8��]Cy�
@,���ٍ��~E�b^���+cϟW�?-���o���b�Nز�������V*aw��ؾ��?,~��ލ�f��~Z�;��|���\�^���~YVw�:Ʋ��oz����܁���R�p���k<�\W��N��
�?���$}gҟC�u'��Ŗ���<��C�hl�`�F
}��p�	��1Maӹ�Jɔ�۾k�;��*	U#ed!�Z�CB��
�Fur��·P7`�[���lI�&�8�{٫p��#($�)vƧr�p4��?a���./�j��u/�7f��_I|^�7���=�����p�c���8U������Jy��Bo��b�6��p�����R���H<��آ��!_�%')�$�Y��%�il��C�>���?����|wU7�U�W-*ն%�Y��ac�B�?y��r��6	Q��Z.;|VU�{8�i+6��("�)�����6;�y�A*�?��8��q��\H�:eZjmI�o\�f6��a���㜝���0O���!�ٌ ���GH$����"�E�l�㾔?A�y�tS�Ռ�]���H0��]H��솢���1����C��0­"�T!k���~L�V�)�|��!c��&x��iQ�2�%�����b1��G㟚�X���@� �8���7��v������!�7��Z�x�qz����C��V$�Ơ|�c4��_��@��r����!� EI*�}�����%p��0�7�[,�չ`��-`D����`����FY-�!�1V�#��1=�Oùtmz���{�������r�B��L�����H׏�(�_��N��v�ҧ"�SD��MN�B�uFJ�^�֎�� ;��{(��B����I����)9Z5/�?j#ъl1��K&*���E��ZH#d��ΣkS�T��(�hiH�aJ����uf��" �s���>���y�A�GIzR�9���<���<X1%��K�<޴5�R��2N#IA��ܗ8<:
@���t��'B9���^�d��˙���ۘH\�Xpk�Fit��jZկ�O�����{���Ma��a"��׀L?@����ގ1R��`�È�=dQ�����iy�+gx��o��Ni��J�4k��s[4H� ����FcW�i�\����I�2\wg�o�"�B��u��<���Z�@���Qܛ��ֺp��Nе	������n�8zt��ԩ��J�P�9R��׵��#�J��J!&#B�J���
�P��ooFۇ;=(F4����f�$�U�<'�f�E^�A���Hpw��a1���P��;ֿ.��S$���v�N��c(��?u�z�)�S����QB��s̕�(NU�Dƽ�+�0a��4�� z�0�D-a�|�{���߅eoQ��u��}�q��/jԳ6FfVt� ��ަ��$:sSbȋU�rl�1�6j��i�L�ZoD�J1t�q��ӝ2�<��	��yh�zx�$������|���ft����ݽRmZ��Zx��������h!Κ�w�5'do� �1:@�����?��ųA������'�H'��O������YB�_a�BTM�3`�Dl��o����4��}�jvg����+VAeB)Uox���"��^�9����������T��ɲ�9�ä��Ś���ֹ��1�B��E93��b�cGӋ�^��u\��ſ䣶uS���*?�[:_�/PP��r��Ij�#�x\��bwŭ�� �I&09���]��#�{��T������E���Y[�Rŷn�e�0T�nuDk�b�w�E���-c	���nfk�.f�D ��'۩`����)�['\[+�$1ݤROP=�����ιK@�k&�)�� �p�$��"�ZzI�6#����l]&��=���a���������1��9R��Ѕ���
@աf�ud��[A��P��)?(o���b�������i�W�K��E9����3p�\}܀
��P*f��K���`ܷ����]�#�����x��P~|Ï���-�Pq�����9y)����)��A�]Kݮ���ͬ�B��(	��?_0=%iL�Nf��9f�W�v{�sQ������u%�+�s*��S���	��Zv������X�P�X	�Q�O��?�r��U���(��'۔��7��D�m���%q��vN��}M7�y�No\�~qk���Y`��s
�"o|w�j6�k����f��9��O�Qo�x��a��sO\ư�x�2/h��TW(=����gp_�W!u��En��-�n���b�����j�����d!��b����&�=�	*kÑ�)r�C=���kV/D4�g�~HI-Q���";�a���8�������+)�,�v x�m�ѓL�r��Lʴ��e{��^��*�
�x����2�Ò
��˓3L]�^����é����R�-!t��n4@E�JWJ�KJ8A^�,*�\��a�X*	~��2:�N��� fan�G�Y�<����M%�)���1��V�
3������.8��|ƣ}
�-D鄵��¶�I�_+l$�m�#̦6�t�)y̾w�n�`�^~Wzē�
���ꍿ M.-�hr��]�/���z0�����[_�@�v5�Q�B����'���4��w輨_^!'i�6U�X�<�\L��{�c��@|b�|{nap�h��7�o���υ�<��Di�zGU֌���O',?Xӭ�]��o�?g�=k�����[.H�łd㊅a%7�$%� ����������=o#�6���f����<�֪I���, ?~ZN �&��Z�'��϶���Y��q�c�gj��r�LZ���#F���>�,i�?N�Rؖ�V3\��l�8RNW{�3T�ժk��浰q�/���{�dz�G�P0W̪�7Q�a="�l&%\r�ǈ�)t�,�����ڏ[8ũ?���L��fћ��O%�|��5X[�yY�c@�ω#h�H�ViI6��	gTf��T��K�.� d�uD�/AӦ�|�\4������Y�B��H_�7��@֐�*�n�������{�f�Y��������>��Mq��(���C2�=7z�5\{�ڷ�^�1N:�҆���r��Y���g�3MooLU�٬��
�>�7��;߲��/�c��S��"��Ģs1mTH����8&�u[!���Y�79�sI���W?D�϶o�
QMv!����O�e�pX�r
��?5$�c=e�$"�mXĔ``t.�h���e�$�̉��xL��hT������7��e�rwd���e�!�a�e���[�22�;G�E�\9�j�H�� �Y!�#�X�ǈn�{�)J��>My9��a��9&��c���w�������B4���Kg�F���<�t�P�pK�{�X���0Ho<������s{�uS��V���/�Q�u#Ke���	1��Zi�=��h�%�89=�lG�%4ʐmk0>���7�V��ý�����;S�Ԓd'{F탈���	�<��&��M�C0��.4�~�ñ�3[H2]�\>����$�'�di��8����Is�� ��͑�A�����f�ꨌ�ECYb\?�ȹ6P��[��8�gJ� e����h�)%D�֌����T�%�9*���\���'�QWR�����7�#��7Y�V�A�W?J��=��3�C�9K���7C�h�sP~鈙�ǉ�E�I� ��U� 0��n�1�pBFf�LW��x�1�d���?�M�	"���{��<���gb�� ��t�"&N<�QRD�%�f�����ڻ���m��uc\u�ח��d�oȶ��w5�}&��d}k�*��g�z)MXp�hh���D��0�^����S�n�]z�,�@����т9<}s�<��T�s����t�<*l��ݜ"J�SK]Ux�}�'�A�(b�*������+�aBZ����/ ��xp9�$�k,ٲ�%�c'�ோ���}��y��I@�d1+	 �o)�f���G�@/�JK���7r����!�4L�Ò���������;6]�'��a�=3��G���%V׷/�)�B��l���hL��s���
	D��'C��I7�o�ށ�%�:�~ܵ��U=%����$JU'/V��KS�N*0��02�D�1�|�s7>������$�D��_�?+���ǈ3���m/G�3�  ��IU��BS{o�0�p�VM��M����ۯ�P0���)*�ZN�vvM��i�Dǟ�GP�N4!��`Nc�3�|��M�LS��g,Z������BN:1ӗ4ZV���N1���~����챡0����hI
籥-.�\/�e�S�����Z��M����)+ٞk
-�a�Y�u��mH�㪚�=�|�UH^������O�ts���2�oPkF�r�-�c�Bb?�a��6˖J�L��UR,	��~=$�9}�*j2��l² HB9(#b�0���t�7�J4�"�Pe���ߚ[�S�g4��5�-�����$�!�W<Q<��@0��8�K�t-�oq�P*�0b���e�~��ݸ��P�?���� ��EZ��h:)~N}���� �uզQmK����c���6�7�=1�BfJd�C��jU�~�loc�	�s�2�ݞ��>Xʞ� T� %|�M�6"�(�I|<�op��.`A
�>��W�9����:�i�u�����k����2Y����������o0�����|����G���J]񝲀�z�T)�Vp������˿z{M��w�'툵���K�\�&�$��@�
�!��bi�8tF7C�(y�e��z��4�w�_t��!񑰸���7k��m�xq�K�ߋQ�bS��T����ɠ���^���m�S4�Iը^� �Q���n/?��5����Ia�����*�;UN�(����a['?�o:|,�^Ũ��GI�(j?R������ �Xre����<'��V�*�� ��=�zD5w�%C�|7!��R���"��]�R;��`5p��L�^���,Oo�A�����/��wN�*��g��lCƗ
�<�I�HUb/"�h�oipz?�k���C����f
�y��g�T�9}
�3T]!7���L=�$(�o=z��>N��-:7�~�6�6Ա$�4�f;nd.���>\�^�z��.�S����t]����em�Z�2�h4+�J������L�J�$gNS"��22ߋ�1r1Z���>g+�1��6�K�~�������D�q߇8���j���`� ���14i"���x��
�K�����@k-����z���
<�J9|����A���ݘR���j	��H���ﻌ�0P����h�Z��ۙA=���3V' w�X�A���	�f�;���Zr��	?�%�~<�K3�6-�,U�^���[�P�b��Є�Xw�y��b�dS�lc��m�q��ld�>���%zr�b�@�8���c��V�'99�`�<�Xq��r27��=�$��6�r�;���K�/�0�� ��Gp��s8f���*�>^f�����a�cQ�l!��oP�;܂�{G�r�/LCհn��a���t4�!?@/K��z�S?�cQycQ����#��ivƅ�f��>�.�
G�(�2䒺�de"k�E���]t���c-�l�[�s��k�S��=�aC�gt�:��f����[�E��T樬�@Ọ�S��z��'�W.�>�e���ϚA�+�º�>n�w�ؔ���-H2�P°H蝏�heS:�s]��j���+�%{`��r��VSV�=?��b����_|�4D�o�	8�zS�ؼ��y;~�?p����.�����.a���ž�3��j���Jݛ	4A�A�5@x������c�>�Ո5�fa�|T��ĵ�N�3�~���7Ruk�_B�6�1�U$�&S����,�	2ϱ�脩��~�b9V0���/��ߐV�)V�q%- Ra�u���U��ou��EP�A������|�Zu4V�ۚ��A�Қ��ճ�Ar�����UR� ����/wF����}%�7�ˁ�c��Px�f�02<0F	���~CJ���G��C��cf�v��mR�����\{��a�);�$���_,�Nj��s>���~�	�)t��mAx�D��{��Tcb�|c/Ïd^�Β��I�������,z9���3Y�^si�wb=�S�*&��G*P�~NYL�C�P�]�{�P�f�-�/nJ�]2j~@��$������ ��L�zPY� ���06V��pM��� �U�9�(��H{���"X�VS�X�����)�;s���"%�a�ڨv#x�UJMD�J�B�;���g����N�tjC�d5�[�V��6��ٵ��3�r>$� ��D��^�J.��K\�����
�JR{�#,�~��F3��Ć��S(Z��"���p�Ѩ ՟lR����'��::�vҊ| ��n*�oʡ �#�#P�[G���� �!͈B8����S�_�!���;���"��������>���1�&��Y1��\���s�k�6bR�n�u�sV����/'����ZQ��{�#�Sg"v�I	�TX]�~1���|~y��l���B�u�;��s|�������G�1K!�Ne��ո֠~�Tj�j[�0��K�L� ���i���$|�P9SY.2İ�W��K����z��2*��;�"��W�	��N���Nvиv5��'��5��5#���/��u��R�rNs��ȡ����"G����uU��Fb�(U�"kl�Bl���5bVoV1��U���js!��f0�U4`1��7/f��9�G%�.�8��0�����'��Y��)�#��bʂ��9k�V@ZFO�mJ��8Dd3ڶ����8�e�b�� �x���t�13/��9/x�u0m\�@�i�D
�CՁhD������"�`���?�aW��mK{�ĸ�8�u�Q�h�7���o���L���%���2��ɗ���hڀ���Q�FVUK�D�W�Bp�I�Ԕ�O�n���5�p�T��������w*�������.�
���,>�q�Mv�x��F�0��K�>�m��qc�k��T�l��QT}���o���mr��Ef��WN�錷[�Z�R����*��*���8���N���B�"�T�Q�b�)Ȩ�!C`�嗔X�)VK���0�4��y�r����W�{v+��yCMx9��	�){|o:���K���y$��F�`��$������Ǟ�eWN���~T�P����)���t9�n�;R����q���4᪪��%I��?M�=Y>�f�}�E����V�����Ca-+��p_�:]�QX�R;FY����!�8R�*�{�(�-�F����̂��9k��g�sf�+q��"��L!�(PQ\o(7TP��'��9��N5(,!�:̎U�[���1�Z�� L3��-��ӻ9i��?*;�h��D܁br�L�݀���&{W3���r?+��W�s��7
�%|�;���B����cF�餛�l�J�����X�x`��#^�.P�Gi��\/&v|�!�C��#o�m���/���p��C1��ي�[T���(��@+|t}�⯸��qV{�Dtڃr��jڰ�k�^Q�;��<�ڃ't�Y�J�C@�_���|>����&����b�������w�K�w=��#�)>���{V�ac���oGj�mA���B�oAŒ�A�ϟ�kg9ѯ�9x���%���i�#rw��v�̬�SB�-���,\�z/]��D�:����=��^��'c*���p.*:��B��_V TT��Ǹ���s�ى|C�c�]
�h?�~�tQ4x�(&�EԽ��:��A����1���%t~AKj��6+f��M	��i��$���CdE�<�Wj��d?�R:��j�����k�����i�Ӊm��5�Y�6g�ӕOnH&Ny�a*H��E���s%����W�D��{W2D��Vx�=�;�8V�����;� ��Wl�6�܁_o�Dd�͢�;ne��:�	 ��2�o$��|�&��E9�n��"�=
M��T����U}�\Z`� �^�(ǥ���� <e�+r�p�
� Y��6"{�"o�'�Z���v���5(O��6�\F��(���1-��r��j�uyʈ=�����P�Li>u3-r�����c �+T�q1Z�����.�/'昿��&N��s��,�A��JJ���I� NN$M�ߧ@�q���G`,awR$k �)�r��	��	�CO����Z�㱣����C/�������'� ]��A�¶&����%����Y�� ��qv����3e���%���#7��Ib��R�SS!�_���q��Rk���g"9s�^;7q��h���FĿ�\v��5�h����Xe5�r'̢M���D��2}s�}%f����g�õH�Z��bbv`��-Y����Rp��6���`�]�z�v�gXQ�jL��VC�"�P���l���,�B�v�D5G�D��D^�ʅs=���ة�͞��l�B�0H�EU��^��zm2޿��\ջ���߇�����'���_�-�3)��g�}s`�Z��R�j�>��-�{>���	�#w�YC�Ճ��k�.�(};��4���Q�dl1u�ѝ��xx��uO��[����"@��~Vk�Dj�l �IQDcS��u$]k�L���� f�
u�2Z�1�B�tI���	��ܫ�6�B��������9�vB0���@�m�\f鑕�n��/53p .I˽Ѥ0pb��f R![�i�UG�xtޠ���"Qt���o�i��'2�����^�~�H����\��z� ̏�վ�i�
P���:�>��we��p ATgM=<1��״A���r��KZE�x��p8�.c��C簒�ݒD��kAbt�~b���
�Z�i^g�����Ut�t�E��)g��&Qu�0���whr�{G�Z7^ĆK��Q��'Mq�q;qv�$���8{G���9U��$��i����UTϐ��$}����
HfdE.�'�L�I>��7/6	DO�Ј�#�t�x��!
�!kz���f�7G����L9ctf��M�p�֓Nj��Hm��/{$J/�b�2V�����J[�ޙ�C�&EBRX)7����{�}�+��\�`�rfx�r���bT�>�,ʁ����c�q @C�[����$W�	�T�u��C\?�<}b�xc��u(>��*f������]���O]�ԩ���c*�Pe�v��t%f�H.x�05�Vȱ����89e�� "_�$g��+?G,;��
g��L������wS�x���-��%A��>���,��N���Oh�Cn�q'����u�pY	�r;�x;ٙ���h��ܻ�������ł�uf?��bx jZ� s~����ט�W�t��1Hm��	���4�%��Ѝ���@kƕ���.���X��z ��S w�/�D���.�?�Oә&)v(�����X:�CgX�@�X|̇�Q�kF��pU�b�n`J�MP��jA��[��e�B�;�ӵ4p��Գ�0�8��f��^O8'魭M/�G��^��+x�Ӑ�=�k�FZe6�P5�j����"����Q$��!Q��a/�b�GǠ�������\��9a!�����FG���{����t���b9�6����s�זe(���[�|#-��o�ͨ�0ϳ
�Dh�7c%���~�[�;� C(��v<+�}T�bbY��Tk�
5?��(jx�~y���Բ~���__,�;�q�j�5���c�O�)S�2h��ǥ׻�x@���<���B���"i�%�v�;�Ar�����ٰ��'��>�e�~�ۯ"�̒P ��V�����ɬ4���{T-X����+D��勏wXx򳰳bй1��z�=�z�r�#�l�_{����%�}ʬM����ĺj�M׉��P%\\�,{��J���gO��L7_g�!��;�.�8+���4%�35��S�[r��d\�|�Ԃ��~��
Y�U�����A�l���j��.>�;_f!sS�k
 �
�v�7�7�*[2�V���v�wՇ濎����E��b+=<>�����qn��+��*D��Ɵb�ZH̥�p��|��i^5����~�ȟTUrǜ�n
�>5��(�tb};�y^d�~>3M(?�������Vj�E�|��_xK# Q�nN����IV5���(f�����6+��c\���H�Ԡ�X��i��� [��jbx<�5���.���9��æ�h�;v�j�%?�zɲ�i�%��v����ƍ�t��s0ځ@NIL3��nB}��t�2�_eO��y�a����<t7P�d濦bv�6a͊�݌�|T�9_W�c��F�!�m�4����eH�0�{Ea�N���4�{�^�9�bo��/W�UbM�q@� c�D���T�:����[��$}�
n���H�B��
6��<@�϶/It-*B�Bq/�^��n���QV����`�Թ�c�"���=~Ԍ�	q�z�v�Mu)���ą+�8M��[M8r5����PA�fa�hs���eQ(WF��V�����\
�'����~�~ە91Cw�J������Y�ci��r^$f��|*���R�sǸK�Dk�ó�*�h�i:0��IVx��<�J�����1��Ľ�\g%�E�,G�l�\���J�������K��a��!�@����d>_� �Z��m���v:��.l�9�S�����pc��/���g�*@"������"J���d��Ė��":�$��
~�K�ca� �i�g\UҔ�y7Q �Nr5��Q{���*+�Ⅲ!�K~�Y_ѕ�g����rضyH8(x!�i���(��X�@S3p�'s�$rX�p+���ཀྵ�m��-0�}�����|G�w����L&�^��v����Q�0�2��#�jx�3F�I���W=l��!�YGv��󐤣(ݸ��ed��M}���6�\���G�2L|�1�� *�7$����a:2�����ɏ`����o��P�]�IE��uS��Az�Gf�#���29ڢ�)�
��A��b��.L؟�m�2��
�l��q,��{<7��{j�qb��FH�F�7 �	�Y�d#�\,��5Oٞf!��]QR�#Bb�,N�-tǙ�pN���k;n�Jg��@E�|�ٹw�`����;诐*-�'�	DUS�t �7����3��z��8�U�!a�  �MF���ֶ��/�H�:�	^c�����(����߄��E2�-������Vƪ?[أc)����mI�~� ���& =�V�ӕ��h�_)�p	{���ZHd�tWL�������Ę�܋�_r8v_Ȑ!jM��I�����rayJGX�r)+�t�2�8���1=��ӟ��tU�����f�e�y(�lY������)c�=���J�&��4���ԑm�F�Т�k6�\~��9rŖU�x5�i�v=����7"!��-�U#�S�Fe������Q�\�O���<`�������1cv���@� �aj̿��LyO"5��8�Y�b���8�G��ӧ��\�hx�&;�o���1kH�x�XDE#d���fw����S�*TN��yΓ�H	�ݥ}:	+5vN~Wz��L+�>�kl ��%__�ID7�
;5��/�>j�s�1��u\��B��?H�ۖ�fK��T��?,]?zK]���+������<c�������b�UA����᱇��2��v�h�R~�.0�h?.T%���U�2KA�:Th�a�q�V�5�[���r��Ѫ�� 't��Ry�؜i�Wd�lsf��0~�z�eI�T�dS��˘d��1�=l�����b\���x�&ðbg�����@
r T�`{����ꜪM+h�-\">o�=$��)�6�ֲ`�����쑟��g*�g��Ӏ�uJ[�w�A�*��X�rۚ�k|��__e�&��8
{)�WSgO	�?��� /MQ��X��J�#���k�Uu�[+a��^�U�o����ǸhWzciȣ����R�� ��NԆ�F}�jD[���^w؍J��cL q�f�5[��k���S~�<gLw�	b}f�
5�u��b�0A���${�g�S@*6�U���Q�����Hzu�]�N��ܾ��]x�/�vd�_̼z��Q��ڌ�[�qbೡXs�V�����d}A,5��F����r��Z)F�5	d1�16�ƯI6v���!� �����=7Aj*�r%[z(ʈ�&"r�Q㬌0�7���_C�����U�"�ˎݠ��9^�"��E3`t��f�o���b�����P�LI��K*F�h��o9�)Ê��,ş]����R�U��31��?:2����:cU�I�G�aNQ���BY���Xa{�	]:c�S���9.�pj�b���5@t�%�t�!�������ж `g�󺼮�(����z�=6e�� &��p`��ا�RԐK���\즜kFv��[��t"�}}������T��:���y����H�f�n4h�e�\��'R{���8c����t�b�{��o"b�1Nl� ��1����u�<��p��~�0�d1�/t� x�]diB�77p|Q��L���ݷ������Lu)*v	$F�y��k�]�[b:%J3����efn��^k����f�������$�R'�@�@u�h̿ g��N�(Z���;�/��#�_�|ǱSRmT���u��Y+��{2}�*���$͇�}��cao�+��ņ�f�%��
�U7�<�VϞ�����s΃��ވ�\���VB���t$䫋S(��"�%y��6%_�Q(w>�眛6X��|�:ɇ�M-7��n�my��ev����9h��6��&�ZJS��BgW�Z)Ҥ�~�#`��!�y�Hn�!���e�\��Ei��E��Gr��u	��2r��$��`\f���!�����
�dRZl�#O˷;�sO�����Bo��Z�5�Ϯ�r�/�2@h��6����,�Ԯ�2R��(��D����c������N�.e��xm�x���t�
�={�{[?�4{Ib>�q�yQ�"I�d���`Qv�u���!�E�H�KV,��`�<��������R�z�����g���� ��?tTM�'�I�;:��8�3k�q�]o��ٷBr�5�؂Ou����)quL��8#�����n?�����a��׎ϋ�����9g�W��=���� d0�cj�)�(�Dc��gD\�z߹�O��I+�\�����f��$1|y7��UG�g_�P����/(�I��l�|F�_|<���������N�	�GZ����m��n{#�TɞsW�/.~�r�
ɘ\5� �����=�nbw?��P8���K_8��s~Ӧ��9�Byjcvf{�8�tHD��}��2s����J鯙ÿ'�?ɞ�&w��Pe$�+�V*tD ��$j0��D�8���|��l��{������ǱgH{鿠d$*�_���ȱ)@o�Z�js��(Qn8�O�1ξ��ŧ�"�t��j�<�D�lA��~����jØ%�Y]�`9�"��1���H_�M�I�P>��KЪ�{�
�&�a)���<6$�J��q\U��� �B��]�|y����S��
7{U�ϘM���{e��5��əNZ�i�_j�p���g�qL��������n��큶pSA#{\�'�����%)WD�	�x����2f��h~K(��D��%�~�})k4SGSv��}}�'��8��;�@"]�(�t�b�p.�x]����x.e.�B��?59���1v�s��rA��x��.��9F���t���	�Z�L��:c�8�:<��ޠ8�0����q&�I'��]����=�Btd�<
B��oذ�����}�;�v�U�bMX�æ����[���WZ�J�;T�+������\&��������,a>�V<�p���>Nɋ�?C���Q(R��[Ѻ�[<����L5	J¼�Z������28OT1�%�����Q.=�� ����L8�uҥ
D�Fv�H;jq|/�b+�g;�2�G#��i]��`��+~�{b��8��61+`~�ݰ�1 ��I0|!��.3{������x�0����<٦�]t���4���o�+f��N����0kc��s��Gw�m�H��zIyk���x0��3����x�+F��|g|���}5oP%Zo �!���3����5,�]���M=��7=c�x��5`�Kz iQҽdXF��Tnp�u����yg�mV*x�3v��k�����G�v$c�5���;�wc�:�ު#�a��p��^{�d����y$�3�P8>}Dߴ'2
��'�d� 
�:�����ئ��Vbjr�8ΞU���(���HA2h	�Y�<�dS���a�����Y,� g�̯S#��*Ģ�+qV$q���
R2�]�!������ϳ������,�l�z����R�+(��O�tV����؁�A����Jh�8�~-��h��BC�+3�&]Pbr�"��]2~�p�@�wﻋ��uhz�G� �}��4 ��YlH?�h�C��;2%��))mi�k'dh�nZe�a5���e�F��W�H=����D����Ý�x�b�,Od��p$��no��>sn6��ZuIp�r�[�Ǚxx�#� �������U���L0�,���x�X�������{����H��k\���3'6z��e�-K��z�j۾�v��8�6�=�^�`X�'���#wL��9<i2|�t
aN����U�l�	-��}x|�^�ug7h ��Q���?f����G/��
Y�l�s�������R=�."�	' �`�<�PͿ|3j������5ϔ�����<��f��Np�R�)��	��^�E��c����9��F�~����� ���{��"��XD>i�8 ��ݪ̼>u:� K�:��>Q*��Dd���7؜��7���"�w}�}���[�,�]��Q�߀�]�0T�l�.W=t��4~ �t���CvZ!î�q�5pL~���p�1��{�E�n>w3��]�cz�*��&��_Pm�AU��LT�D����>����J�u$�Ow�.)x'�u�ќ���
	����I=ߝ���ى�~��Olv�X���#����Q�Μ���\�>����;�i��,t�qB4�
mm-N�7P"��9�Lp�_?�!��� �zt��ڍ-/]uߏ`x���%�ة�ɷ&��h��Z��U�I_P)�^�0����6����H/��8c�Y��xU�TB[����8zA�4�/�8j/ԋ���S\�2�ee�g�T .����=�����|pa�"�B�2W]�����~no��Z�)���M"��=)Et5G�/i�.�6����嶺�C|yWS�S�����No_}�����ߐ˹Z��� 8�1����o#�%2��	0��p��6^�h���S0c��~`���3�a���襰��\�nS�u���%��;ǻq���E1ǌ�"$mNa�!���M���1dZ7\��z��(l���O$�[�Y���f2�f��{�!��Z;�"F�R�hg1�����m��_`��M!�,�ZU?�%@�q�'*u9���^a�6+���O�0�
�B̥0��r�O��O�!�BX;v���,a1��0��r`���X`�!�R9G&Dm\ۨ3�ׅ��i�xצyS�w_�K�5u!��?�����6�f�ȼ�Y�Z�g��GL�����}�����H�6�+۽ꚝK������Yˡ��L��܆�kK��8N ���@�\u�z1��&/,��4�+� �][!��Bq�P��ނ����]W�d��c�g��c�U�e����f�ߠ@�l �h,Ԅ����s��*�iE����K��?�d���q-A�}8�Ǎv� ���p��O~l�o]|w����@���`L�F�6����8�@�fs|�꿕EqӍk�[�>umh�k�~�H!s�vM�i�9S�����F�O? �\
Z���l�Ѵ��3ݕ���˨��!�%�QRJ`ҍ�� ��W�)-x����`��D�C�'c�J�-���%�3�u&�����%ϳt.�]i�G��~�V���}��8�����mk�)S��.G����6�1z*���I]�d� e���%��pX�7p�/ֿ�sZ��D��s�-���t�vT{eE����<�n��8���fU�?�u^ZH�e��W�^к>߯���R�2	~F�q�1�	4��B�@�.�񿢰���;�ZKl���M��/r��W�zvmP����A|��(���A��m���-t��@�ʇp�.o�t+�J-ԭ�u�(iu���Y���	����I�Y`V	�f9+�Ob�Yc ���Z�����S�t�����ζut��
�£ �!.,^�G)v��uB�Rd�ʟ�;�^��/x7'��fV�'V�/�Y騗'!��(��,	q�����3:4�}����p��{\!�����P���Rz�5yf�5�o�:���=��a��]�Mt��K�YԠ��VLp�8�b��t�����k��z����:,mqC��0CZ�/š\�Lݖ�ѾY�-ip�����}݅p��"=��O�[hZ�7�+盡-[ڀ�Ћ8 ���]�G�*CX&��-��L�5+��|W��{s#4��C[�@&��8[ �I�R�wc)�� g{�n���<m��s[����ۓ�ځ���4_P�X!��n������o�,�U�s�RE���@�&V��᧠���|�}�s�y�}b��-(���ۯI<�H���Ni���W����#kSX"3S�&$�;�Xߋ,�)��	��-L4�X"���A��zX�J�ǹ��$����(]xB9H�Z���@��P9��ai!�W|�=*�r*�z�D�_�dK�e�M�N�S
Kly��G���C�s�Q=��2/�o�Z(��GtC7r��~/.<]��I���.YMФe܀��O�3��}�(R�Ѫ(��E~J�v�&���u�m�O����a	�t���ߎ��:�<�n��Cx�o%�͌��Pr�d�t#\�"��6`�-w��	T���	4�Ǜ+��:�<�;�K) MΤϟ���)jM�Q.p�ZR� ��h�lEJ���W�i<����f٭G�U|�u�l�:L������z�*�]�(>
�5!PD'/�����F�C$'۲quv�w�鶙)ѵ�[��ad��y��]��J���s��^�9���%�Yq��K1@���
Úyy: ����J��~zq(�q��/ZwY0�4T�@晛�1���� �{s�˶����q?~�Z�W!+�*@�v�l��DA�u�R��lz��:����k���N���	��� �]�Z�8��{��b���Un
��FH�Vy��>}g�:���8�>.n��F�Be�RTD���ugS�]t_͟GY��ZB���U.����eR�4�Ϸ�+ݭQ��T��벩5��g�d:�*
M߇�����l) �C�<!� ��tZff�5�kgC-��
^�.������= � Hj+�PUpo�D��� ��t�@�=�c���U��|!l7vm�*y/QȢ� �:�T�{0֦g���L0�M��2�%�ď�l�,ӧ��$�qH��6��{8v�����~L�MA�M°_.E��P:K�t��:�n_
�֯f25�~�<�^b22�qB8{���E���U�9eHd���s u��L�#�@�0�O�\x�Z�Pl�]�[�QH���bW�Ihn���ρ��;,A���8��[����������-��ip*_�9@��y+������`"�w�Z���T;� v�8TѸI?���f���׽<~O��ʷ(i: ���j�b\�yq!WD�R �'�L�~{�&X���� J�cb�B��*��63ڊj��K��R�� .�]�*�n�h#`��ƀ|�2�j��;���O�g" 	{��Od��\�b�;�Z�"�>�`�C�y��*_*�^�?Akһ����{$��I���ƣ��U����ݣk�n)Q��ڭ,�:s�L&4�W��_V�h��m������,P��s!�6g�ҧb*��U��i��� �V����71$ %�-{������Ѯ�)�=>�;��9=n*a�NY����'⫹�ry\$�_�  9�C�Ďg�\���z�\�;�*�E>���
.��Qe�v��ަ�A�tw6���(tW���$L^���"�J(��Q��%y�݈����&W_.�u��Z�&��Z}��,�jI!U�B��!Z��`;	V[���l���m9�a�Re���~#��va�}m{X�Oz�;�K�uV01̿��MyS�xk�&�d�V��aGt�� ��H�۾H?�n'vx�)w8j����t���l�~W1S/��9lD7��D ��^n�][ر~՛7����_����}�s�J�E�@P���ҏ�a�!�ܔt_>U?���S���&�[yP����B�
D�.ћ���#�p�&o�uN7�`�w>�V�b!�c��I�{/���9Ě�w�U�����
C������o��h�;8���e�$���k4k�ua�+���mS�J�2�=Ɣ�@�4i�.E}�u(��MT) �����ͷF�yᰓ�l¼��z�}�o�Eȸ��3�w�[-q%�I�G2%����!K�.�c�F곉h{��GH��2�A�]B�e������! �MN+�
@	�˰�dm���A-��5���9wЎ�����f%�
��E�{!�H-���K����b����Li9�� A��TCu\֨�v����Z�^�hs���z��{c���~�s�>���q����yrLK�/&��IVz��
j��F���Xp���C���4RK�?W���'|{+�'韢�<���j{k�5���a����o���A��#�*��2��k�C+���iX��L�q���)2>D�6�yD����4�b�%b�b��:��Z& 'h����������Rn@C�CyP=<���<�k�pT<���vЏH�K�����F
O�Q�����[Jw�g�P�� �f�ǅ7ރ�j�C��/l�L�a��΢����
����l��FTC��,����^X
��[�1���<��6�$��@�E=��m��x�]�l���)��}#o]��VmCԨ��P tB���o�I޺���������]ڦ���r�L�A9!�C�a�=~�8L)���]�y���OQ����Hʷ��VzE]��S�~�[��8&<���v�w�[�H��Oо��G�<#\��'�-�)D��l��i�b��@�p6s�$y����ȉMD����j���G_Pt)�d<5�������B�(5_�; ��v"�6�o<)OP�a���TmwO���0#s)M_������(-{x��{1��R�G�U��;tS���\=Z��\�,~OZ7#�,Ew,8ԍ�j9ᔉj�YW�^b��.�1������FQHZ�@�r� rԉ�Ks�����ͥJ��$�4�	r���$��o��S^�N��ռP� ��!Y6��0D;��té�KN�;˧D��]%��gdtH滂H���?����� ��5�G��<��A��ϑ|����Hl� ��{��$ƒ.cv$߶�0[#o�A�3���V�����"�Z�?�¥�cfw�.{�I �	(r��l�w5�>�^��s~��S�uI����YD2*};?�N�c�HR�GD&�ЈS��C�z	Z��3��2#�S�,D�r8���qJ^�4ŞUJ����ҿb��G���n������F,� '*�,2gE�+�wC��)�f��'X�ӂa����˱�7́#�$ؕq ���|Ɔ���/Sy�qϛ���ʔ�W�&�-��ϩ��������tK���'B��9�YAፘs5����Vu!r7'F)=��,�A&�?f��c�lvr�,�3���`NBKDD*qE��Wvx���Zbgv��*��+�][=�(�rh���,����S���$$�n�jA^�кۓ���Xa���/�
�f� ���2�H�ARp���c��w���F눼�ʍ��8�aU�(���}��4��D��Ǡ�e!�	���乴�N�J��<���id�0}�z邮�fn5�Q�	�����抡h	��ieưC*��F��Zd�b�ʸU9�+�C���n��?"Q��FL�e>~�����,ð�]�kb�z�7N��T�$^�vيcw1	��B�H9�� �M=&N��!M�O�O��m����wJA��os*�x������kA?�`�e Jly*��$��[{�$�E�K1c4F���>�@�-���I���Ͷ��Tv@�V}�w�PI�Ԓ�^+�Pg?mԽ���?:�C��-u�nAT��9��ڋ�2}����b�����9��D9��u�b��73Z&�VD�J�[hX���x��`�N� �J���8����J1�V_��v>�:e�L�����m��I�Έ/�j)*K~+�<��T�?��b��Y,ÓЂrv�$M8���Aý��|�W�刽��6�(}�_�"�F���`_�؄�6z�+�X�	0V�ee<wq�������s��H1�i��K��;���
ܙa7�~�u߿Ȳyz�g��[3��~/�?il��˛#�����]#�~*L�C+�i��W��T�xu�=,rx��_������w#H��x&�,��F�r;�]�8Jϩ6Ȯ?�n� ��HKOS��}���S��)�v1g1%_J}����2X�%��)v��,�n��MsKC�*S݅���z�� L�5�(8��:'�8�m!&t���!jɯje�S�`c"�Ӥ�t��P�PYz�H-`I�|����@�Q�A�4�����|u�#,�W?�#��lň��%�y����bѝ�x��k@�6�K�J��G��f��L�R����|	����(��|�ۓ�Y�I��ڧN��ω�����{_�l�t*�'����$�U?"{��_�y3HYw�B��m��G�:0�W�^t�S�O_�
����K�w���n���a8y����1��c�tT�ឃ�����.^��c�I�l`�~��~`'Q��[2�!�[I��bԻ)��ʓ��*���W��@H�S	D��e�Ӎ��g���u=�rX��e�u�镄�a��E�δ���x@����d_����,u��:��rj�>V>?J�#ֶ(�������
��Y9 �G1ҺO��I.|�(������s|�お�Q���^?�=G�]e핳��C��gP
��w��9��r��U�'
<���5r7�I�FXk�����j�>I�|}�V����ᒪ���Hu��׮��cM����M���Q�x�F'Ip
v��9�v6����l-�Eg�3�@i�<��VQw�/J��B���a���S�]�:�pa�5f���d�;��r7������@�����&�j�}n��M"m>����aL�,�{�7d����5�����>�p5n�k۸@_C��9e��~�2X�0.�����(U� �-
��e����w�?�v�&{)�dk�!�pC3�]�(D�x���鮼�Ņ*J�t�{5�]�F�Wq���d����x4�@����!7��k(t;�w���7�`̝ӥl/E�x�=��V+���My����|��7���*��y�eZYam�������(M�Hj9Hn<�d}��D�G�e����[o�̯-3P,�:ǄA�,��0kd��~����.�r�Mo%)��O�!� �Z�tYWU����+v�I懎�P!��t��b�W� l��GS�RH��n,T�7#�w$��p7B�(� �[�<w���m�kn��Rx>�I5iǷ��eH-]�	�	YH����2<U��w�X�E}/�ݓL�IT=��W�K�V�J��3���獰�s�t��<!�����	)���&�̹+�JN�RD0fо�j��� �n;QIc�H�`$��N�ؓ�^.�Q�'�DJ3�o"��ާ)}N+=����NOl�r��Lq��nM�GM��x �	�[CU�x#��zLgbd6�1��/�����ݸ���X��e{�����oK������_e_{Z�^�1)�� L�dw� 獌Q_Q�OK��8�Fj��4�E㻱�h�Ɣ�I5x��,*d/�#�3sxÕ�!ާ���TK̉��-��:�~J6(�]�S���4�pBOR%��s'ZX�����vݸ�_ ���r��2f�h:�pw?zA�cQk4�D�@w,�UZbLZx�Z;5uH�]��I�sw�ۖ�?W"N�'�ƖD�gy)d01���C��zX�pvմ��ŭ+�IG�Y��ګ�(�!TY�h��G�����!L��=8���M��u݈�1ڏΠ.��~Ķءg�W��	 �s��ʏ�te"	-����uf }�(�W߾Gx�M���������O�,nܜe����	�%z�K:��+<4����<�r�e0�2���Y8+�t=l,��>��$�ql71@k�bF
�tk7˳����Z�A�j�|��L�'>x��e�|����ă#��6yO_ª�ltt�L[�庥���9��uM�����1zNW7�G��6; ��o+��8�K��X;o�=���zՓ�أ���4)l�:�v��~$d;q��|NP�>ݜ��)n�<xPmNx�M��nB:��R5��WGd�|����M�ɬr�G�D�9�']�.�	��&�r<�uDs`��v���"�s@�F3ZF�>`Da\�Z�[���@(��XKd,��[P��"'�1HGe�4P^�����Ȑ�iY����hT�?\�ʴ<O��,P�r � k�?~@����^u��e�@���(��X����K�:�hF�q8	u�{~��<qx���-��6	�����jo�'v�%w���P���|W�33Y���V8����q�҃g-��'l&ǿ��aＲ���@@�P�s8����]�Pj�/�����8��$���N����+'�(V����9=T���7H��K
򍤲��\�|k�FMKr��+4�e�!�r�	�٣���=��nΧ0���OP��Vj��._]1�5G�OX�a�M:^�M�8��b��z�I�1!CA�$$���MʴO�r�2�K��	��@S�n����0`U�d
��X��8�F��ʵ����o�>:�s��e�DuQ���o��Z�u�|�?;b����SC�����V[sY���!�l�Y��A�)z�m�t�ԍ�6� l<��Lt�, =a3j�+�����2ܸB��g�~��H��']<����Z�2(�~N^,J�[�Q�=A[AMRw���}�7X�P#T;�/�8:Հ��?���c���Wu��M<�Z��.<�T/+������}VĮ"rF_��#�`�W��z,}a���?�)��û�)�#�|7�N���B�쎼$_��#�ן��ţ�6�������w�L���R�ҏp!�|��,�|_ ���k �h�H�)���׶��C�,��Hxn�,��ϻ�5&&_��(�RQ��m+k�e�,�+�+m�f�"�������`��� �h�GA�.����Z�#��bR G<l��~!�Oc�f�Ei��o�����y�z&��#�d��i��;���Is�6$��W��<��Y��Eߣ��@�'�JUy�k�`��Ǝ����G���(�C����[_���H������l����t��v�.�#o��@)�w��u�
/R
8947[kf��A �P=���牸X	��8��E����?�$'e]��́G^0�ǉB'���4�W�\QR��?�i,H�Bu_:��Z�����@1��Y>م��mc�S3
����Wnmδ�c�J���U
A� ,��<c�?���>`��o�������p�����K'20�$��,P'w���aw�H�fZ~x�pKXH<Ѽ�=Ƹ�YR<^p�$��S�'�m��[^�bY���k]�������A���;ܕů�#h"Ij�ER��B���/B(B9�h�,��h��<M���j�\1S�=~��l[�*u�ۍ����Q���eK.���u�4?�CʂX�\���D��Z>׉#�	���1���O�݋�H^������ᬑTaQo�{�Q����Č����l�3������Վ>mqʬ��:�|�QM�CC��u��k���kM����αH�ff	[�'nU�z%�A���pj\����cqMlw�����z#�+���ώ�u��_�������]=r]�J�L�T2�v�x�q�������Ԗ��k�6l�4��Z�͋�^�����/IV���[ƃ%G������~����_ʻV���f�4�������庭4�STNu���*�F��QO��C�2H�~�J�p��s���� u<�~��w��,Z���cXL��:'���/��5�WY'!M��N��J)v�w�j6̛s��;V&�9f)
��s'��t[�����J������O�b�E���/�Oy��N���7�8k�c�r�	���[��:�^�n��Vz����uѡq2�?ߣQ0��j���q��_ߝ'��K�ɼe��#7e3|�P)ff��_�ߛ]�����������ko�i��G��%z�l����<I �L�CH���@~_e�w�=k^cn&�p�'1`��A��B�2og�P��Pr�����u �� �E���]�ے�f��e����S���ˏ�����ͤLaT�:���A;�����[<x31:��ч��Ɂ��5h-+H�2W��D��������B3��"�A�/���0���%ɫ�L��۝���-���5���X�(�#�$%�]�&�aw �Ē�x�R�s>?��:#�^�Hu��/��v�#yJ�̏�V�ju��~a�����Cf�@�6�*0�,|=.�7=��g_�8F�ib�W�S�f:����@�A���&;��sǉʸ" �8K��䷺�b�;�]�M���*����[D�2� ��~
}E ǮD���Lt��>m��s޺�{P���X]��M����V(Ag+qWk�@o���u��y�� �c�˜��Y{2�Y��,��@�NP���|�b��(��r.���a��|*��i�~�^	���Y:��KͲ�ݛx'K�tE]Șpa�*r��(mՂ�4�7����NO��	����4�C���T��B�D���>k�����ȗ�FI� �;��	X�ŨZ+:��ɐ%�%*k�@�Ҋ�~���"��=��ˣ�}��ۚ�`�;Ƥ~	N!t��X�Y���a���DgJq����R(Y�C<�>���vۀ��l_���,�� �����<>n߿։wYHvmmЊ3�TÙJ�Z����4V�_����`�hy��t.8�IϠ}�M�BE��_ս���OC�>��[3Ū����(�L�6g�� �/�-�����2�2H���=�s��f���NoI�'�U��p{̲����y�� R��*���(�?�����'1��ퟴ��s���x�?_�E ���vp�(����:��gh(�Ɛ�r�_��&��_��L�)Lf�	B���Lj �<ȼK5�9�'���c�����Z��������T90�5K�ӻx�U���Q�Qޗ�X}�痿	�@}��L�AYj�sS^��f!*�F��ө�4�3�13^�q�Me��kBv��e��ä�V��rWB7��/u��c�r�f�6J�5�s6���૦���������K����%,���Fأb�eZ��{�-Ҹ0����!F[}`��=`��$���w��ͧ�a�������dU��J����4�<���X��7e���ܹ�M��@�Ū ��^�h�U!����͕5�{3��t�gu̊�P��]�:�3�E���Xr�'��f��K��}υ���f�C������A;$�Ӈ`����'���]ѧ�xk�iA_��RmJ���`��*�Q/ڟ����c�|��uԔ3��!�~�nvPIX�A_<!`���A�4���ח��KYp�X8`�u�(_OH���=G�[�W�t�I���9\��^G��>����Y��&��m��PC�L:�N����2/u����S��������ȫ��\�,��>�X�k$V�'�}�Sf�8�v�@X
L��%Mr5��L�4Y��#e��=KwT���D��^2��� ��Cv}IJ�+�`ěP�R��P�� *�Ý3�.YNޥ�0��ď�T��G?o��57��|����=_����3ִv�q���$𸺿f6���=�w7����@Q\Ul�U��a:�^���
��S�bY���ֻ
�"�B���ِ,sG�i�͈y)������.Y2z��f$�$��Ⱦ�{���y�_�a�m&���u
�u;�V��=a�dמ�ԽXR�;�
�B��PHP�.z������X	���Qz<����ȳky� Ő��<*�����|^\�AdKD�g������le���"YP����,O���ᇍ�.�/�pل������ ��+Ef����T	���ILuvj5g������� L�v���
m��\�`�դ�ݝ�%�c��o� 5&�nW�Ch{4j��G����e���x���'�~��fa�-��ƆQ�G
6������ק�dɤ�J�!�]�g�*���0-0�_��Mht��j׹7a�ɕ��,1��h>���^��~PQ 8�w4-�#��c%����+�]�l׬Wh�'d�M��;YS@t�pd�\��4	�ˋ�{.��xK�Cu�K�:��T��̧.F|�y��z%��v�0~�O�R2s��N>�3��e��j���v�U#x�"�É��B\Q�/�u�� gy��/~� ��rtw�!�����9\���-���+PE���<8a�99�9[��� x��4T��Ծ�o��N�H��\i��?�����`dgA���o�������e�:Z"\�癌א>Bu*�9�]� f��s�E0�QZ[Z�+��Y�3n`�Ø|פֿ�E"�$bqw]�+�7�=����vb^����INLL�2���u.n�Fs]���5
5Kԁ�OB����M���c������T4F��	e��{�'m+/�e����x^22��-��>X�G�{��b�[�c|�(��ꐢo>�ޏt�A��c��������M̷�!�+#��i�Y������������g%����DB�{ǭy6Y@HŽ�.7��T����-��%Xh����14>�ͽ�#���V�M�(�����W@�_Ę�ͫ(@�!�6�������w��(N��B$�5<�7���"2�6�˒��i��1��ð��\��lY�ȫ.�&����cs�tq����!�Nu�ċl�,�C>��Ѽ����Ʀ�0�N㸩RϘGoZ�:��M�t������1�d	Q2���L~^�m�lPtl�Pr��x*��IJO}D}����	�&]���|�7$��er��K81���)E���]fw����{���j���Z��U-E�"*�4g���J�Z��j�qf')+�J3/�`V�C:�;�Ng�Q�o�b��clN���nV���<WI
jX���Ҍ��@$�7��:�YF_=�v�K����ئ=�	 �C��w�bq����<*��u�9��߿����^5X�0!�7U��V�a���;Vtגݛ���Ն�.U��bcW��#:����--B^��D�����rr�[�*I�����4OoF,V�pn]�8��hA�ˏ���אJf��P�.��/�1)j��i"�bE��jqİ�liϱi����3��Lu�s4,�.�T�����DBl3>�YY9x̟��ݞ��$ �:Z����?ŉ��齄��]�#P�j4E�D��sK�0���{*�N��υ �H`��^�$�T�󓙝-�f+y7��+�c�v�2��P{r�E�S�<�n�[�-�	�J ���T���$��E�7�mw}l��Д%1Z��I� g�Dy��.L���G�C?���oXW�j��v� V�ңX����b܉3�Q:����	�P��ct:�ݻ����<� ��$9�[�� R��S�=>\�1����?�b�LUE��91�x �MK1�s{b�� ��m�nd ��"����>U-Q�����u>��qyx-��������X��0�%�~��CY���:tO�i@T7�yw�X����~]�㤌�Y�3�O��бaH�^S���6�<z�H.��˶"%�f��=� ���m^	��$C��r�ɩ����K��/��ȵ��<9��.�'�� �X�֒��2�x l���r�B������9���hX,�B%؍$�"�{Z� YRoe��hרJ��c��q������2��l������YQ�*)��0܍�:�q#K��?!�v���|���q��S��y�����~<^�h{G�׋�}��ҭ�##��	��"��WC��3Jc ���&�]ǆ�C���� ����Faܬ�����C<�+I�|�uQ$�ϫ�G�Y�3���x����No��3�b۩�x�����tx:��\ºӔ�2�7
)Ł����ie93�&j����������%��S�A��ȶn�7�|�$���5��t��`�}ψ�	�M�a��/�~��� d���K��� 3R~�z "(œ1+ȫH�vew'?�-� m��;��0̷��4�I������8��ԑ��4𾢬���G]z'�uI�E����(�
zi���� ������ښekƝ�Ր���w5eه:��.�pe��'���D���L�M��T=�Cۋ������"��[\��%p�HU"��Pcv �D�RHV��+�tEQ����J�gG"�QK*М�yll�o2�s �	Y��\˧��,�ۥ%+X�"�¨�kc����ᎇ�������3�G���\�$�M�.��T��w�~��y:����,��Q���w1�q�}]Wغ�z��@��CUvLJ��$��Q1m��
���ị����*Zڀ
��`b�dxK[L�7�c�]*�+�ǈ@��&�+@�sQ��)��-�ں�b&V��`ߘ
�:������}�)4��U�묝�����ߌ$��B8Q��u�t89����=�{�"R��Y@�_:������2li���+#$8�O�D9���z��D����I@���G$U�7Ȓd~�1Bs�����5�l{��j�.r� ���2oBG���3B:����_$Đ�D�i�3�	�w?���fI>G�{IvQ_,���d�`ͻ�7}|o�fI���]2��AL��W�<pl����LioyoCD�5I����*�)���&c��5����~���(MJ��a�6#	J�H7Md��?NU*��n���JA�-'%y1�w^ �J�O����<0�����j��x�B�5����Sr��f��� i!��4����\2���^��������ԭ��ve4ߜ�ƍ$r��#���"��Hʚ��~"�w2�c4��Ȁ� ����5�}�$�9���\�t�M�L-�ͽ.�Y���9�Y��ܩ�4���2kc�Ak2��t韞��0�9)�*����>Ey�H�Y~ �
b����R�ލ�.%X�5&��Ad[*B҇�O�V|�&����
�tqa�1����g�QA�"sܘn�s=1 �Hd
�(E�Yq��w�������u���֜��ǚ����nщ��,��8�������W>va+���,zEROС>;G7��
wK�L�$i����Tv5O�e�GMwڷ��b�"�G��K�6_���j�i38*���/��c!F�x��uQJ�1�u��rl�4u��� �v��o&�ܪ?���
> l]��,ƙT$�u)x:�o�O�&%���¥>�2���E�ȃ�Eɵ?8��1i��x����'27����{����X�! J�b�y�.\���Y�'+���
{Ў>�K@$F��6�Z���"��j�:�Q��"��q�b��H�Xo4
�2��Ѳ' ���seL^�H�__�,[Ϲ��A$	$|�B�9]�~E��d`�c�cs��q1�$�!�n�8��4�w����?�\�/��ć�Rs$�1P_�a����G���B�)<,S�- ��J���AA�B��GH(�
R�Iݾ��D��Oڲ�CDFEoQ,V�@V����ɕ���t9��/�7}��H�/�;d��q.Il��iI���{��j�H9�,�g���.*&$����oO�� �vC�Ь{w��}���n���qUH�cR��ڄ�xsiѧ�ܥ���ظ��ЖS춷\��i��,f�W�t2�;��:pw�N�7d����=Do��P��BY.�y��E��h�l�l^�
j��|���޼��x���$i4��/�M�/�X�؍Ge>��N�D��n�#��M2�x�Y:x�e�t;���#�
��Ì�n��\��Nso��Q��U	#y��)�gq��8��*�4â�I	MW�89�m)-�b=�vv��;�.d�Q���w�z;jR)f�$�~���j��K�; 	9��AJW�Pp�
(����2���N���eP��F,��9(��¥�pp�=D3�q�U?��S�o��Rl
�N���"�So�c�GAƴr��∦=w�E�8����s�oꗨ�[��h$�n^��vfw���mYD[@'�a�;��$��K8�%�t;�I��l>�G�N��
�=�[�0��
@.�$����=����t;��:,o��5���E�^$ �%�W;�KU�Q7ãQ*�\����L�*]����u!gY׷��&ۛ�!�'�e7���m� �{���U��R��*T�\޿V߽S��R�ƥ�:��e��O��-��U孻#m{+�[̋�8��O�~m���֝F�!PZ�.�vK�gMac��A���X�-aD����A�E�N#4K@��?��A�OM6���z�����d��&�nc��@1���p��q�/I�5�*���6����l��pI�_Ț�K��;]��!��	�h|���C0�X�k\]�8%Y��+�š����̐��z��;��G��;"��R:-�����$S��MA{j`�am�2��L�{'�P���CIf4j�A�6��$��Z��+;����
$B���Ǭ��7s1GB8�2P�8fU�GB$*�{�d���)"�#=�Q,����Y��/O3���b�yt�o^x{�R�����@)�(9�A��)M���wY}�Z���z8n\���5�w
���(��A>ɥ�R� ��e@<�Oĭ�)�V�!��q�F⊓��G��u���6����Fm��'=�v��}�ڃ�Q��H�I�I�	N"O�Zn�_�Zͻ�&Kq����s�����@�8s�9�������ۋR�(�_Z|wAc�0y|	�W�D��	�jq���p�L6�v��zn�<IQE߽�V
Z�3$�������3��;�sM/|x�,�44!��,`T��/M�����d�gUR�����(P(�Dr�bu�����G�&@�C�� NNA�,�m~z�ThR�Ӝ���]A�H��ք`J.�@�Pԉ�^&�F|��M��d��]{����7�sl�����O2Y�S�qc|<ݕ�L�\��,y,�8��9f��[,��C5�*�q����C�B����<��b K��?티B��L�&g���*�JXan>�3,2s�2��{�9�g��G�9�|�u�a,&�ת?!Ż=�;5����� L��D�3�@Ը�Z��z�ւ�:�������Q����v�r�!�}�P�f���H�j���֠��MK����s�{+��׾�����՟�ܔKR��y��u6�8j�Z 4�o��Ul��'�!�]X$�m�֙��x��C�^Cnj�G��V��쏒� ��l��#u�0�	Gg!̲�H� ݙ���w9=�Ѧ�%L�A�J�|~@�<��a�._�`�A"����bNJ��&�J2E2nd���'T�a�l4�Q� �2�lC'P�Kx�U�!7'��U��W"I��X�Ȃ���8}x���� 5$���|�9r��L�y��G�lw���%�>���U����+J�f���,�����1CT�^1�����i�N���uI^G��0�p|������ ��]�{!�I{���~$���ED�	�;����iqkFF{�8r�B4�-����8@ih�~ș�ei�oT�AO��Q�0�?J|������E��P�5-D��X�՜..����u�/��A�K���|ç6�G�m�s�A���/-��u*T~G`IZ=E���['�T�VzUb��E���KSVD����!4����{��E�ژ���ġ/���CTU�œ�l�I�򧗠S})�o�{J�$�|q�-�,�ě�g�*Ä�{�O�C,�;�zyҰ�wnyOU�&�����ߤ����^E�������w�3ʑQ����� ri�xJ�@v�:��w��倄+|ނ>���D�֭�Ʃ�a+;k��ե
m=��������L�{D�xosE2Q���{��s�j��V�]Z�B���&���NË��e�����K��*��2�i�`'��Y`Yn[:#AJOv2=P1%K�B���Eq�Nze�* ��-A����.0�����e�~��Eݎ�]�a�7�1S��^������?бS�[�d�v֌��Y?ʻTs�Fg8B�gD���V��2V�|����!��%�p]�me%�NxLv��
�TCM�P۹�����)������1!�˞$��b����+�z0��+cї��wJ���V*�����˞L��K\;�)����g榚�q�9-"�l��6W&<k��aH5��ץ�o�k?!s^�$G�����r��#Q����.ɋ�5Y3]�$��&,��S�g9�,A&�4!d`��vXƾ�46�~��鄃.ğ�U�B|��D5�q�q �¬j׏��U����&���B��r�3�^���~8�.HJNL��-��M��i��`�<F�Y�E5��ï�]y�,�y�f�[����=ňp�W�u��d�����2.gt�c,�ց��;^��>�R�>������.6�ab�A��*i��;�����g��|����"x�9�F��	j$j��B�9;Թ9Γo�����R�)dv��W��M%��Ш��ؕ���,#ȫ�C|��r�G�ɂ��wQNu���nd�9��MB�t��XI|��~�l��^��2;a���H�)�&N�u��H��x �GV�@�Q
�7�;�yI�_�N��aW�X�nW�}7cc[a�MK]\�.���D�KA�|��:}"&m>Ä�g���	�V"%h�n�$�x_
�,p�m�VΚ�	�c�ƋY"�(,�|�]oT�l����/q����"�Ġ��1�������� -ujgX�ڤ�lg��"�Q6h�Q*q�?G5��}�1T�n�뢨Ij��]q���r}��s}qUַ[����� ��R�v
7-Dә�~�������˹���@:���܍�]�X���lC�og������l��D-���ǥ#$$�\����:
u���DL�*���q���I=��Eo��&�j���6�2���o��0��!��@���u��a�W�.Nӫ>"Q���r��,<WX�&[��;�sRX� �Z~P�kQz���� ��Y�wn��_O�C���2��glX��j�F��L�3��"H ��e�f�$��`-JϱF���Q4\���x,9�V5냊m��?�H�&z{ΐ���/-��BH}>$Z��,��`��������~&��k,p#r�%��J��|�=��;_�UI��'�E��D�����bZ	׽�Ժ�V|�U����z;���Ej�h���R��t��Si�`@=(R�ea-�\o i�&_�`Bbk&�P�^���7�W�Ej2p�j�t�hB���T,�G=x/�#��/|i�(�_yJ]��kig����y�s��C����W!A�'U�Qi�6�7�z���jD�hm���M��}�qY����G쌪1t�w�|ǹvl��ʹ�����e]L��7!n�E�cш��M�9����sWz�wHqyi�^\��gs*c{�&)�����8�xk%�q�0Oc^e���Q��	^$	ԛ-��w��2f� ���;�A$V�?�BD(3K���cnO���?�����}�IERºw,�^ǷU�c�VT�� cxM�dN��/.tLǷ�ԉ^V�
5��c��Z�,����G���[�#ǣw� m%���R�*��\������&��I��Om1
N�ЌUeGe!O�f֗���y܇��fm̙�*�0z�V����^Ҟ�$�3$��*��͉�*ux9ߢ	��ۧJ�~��1���d�_�Plb m��aW
�(u�a�g[���g7�x�����	?zd8�
�Tz��!��C�� e�~6W@�	��݀p�`�J�E��>�=k\���kǍ�a����-/��7RRO�R����f�жt�)zP�&A8c�`�֑�ŏ�*ا��]e���ޝ<d5�=���Ͳ��x;�9���"ws#�9�"�A3�j���_8P}�I%GU'~�����#%����V�>tKl��J����T򿤹L�)�_��o��<���hA�E=.��6Ռ�0�9g!�`�Z��`rf>˾o��3�~/8��͒�<�@�ƨ0�_��Ի�B�Ȃٳ����h(��9�K�˟�H_s�b9KOh�<�LpΡ��b�5[[�#�Qr���?�{>!�@�ĢΣ�U9�%t����ۡc�^I��܋�*�#9�8������XUtਏ�������Y�t=�A8�a��ɱ��L���d���p���� �|Dӊ'OCh0�Y���Q�n�n������n���x��˃�?d��ǅ��dEN>�LLr�y��5�D#w-�|� �Gk����\əT^�p�R-[�}~�����y�w��#ˎ��?\�":X� +�SP>�nV����4�G�jw�`��6��K��j��2P#��|	�;�3�T؏�
V�l����m�\��	���?� �
���2&a�mE��+UnA�~vl �K�B�B�b���S���<��H敿����9H	K�����n��;D!T���_����#2�Z���M��/���F>���������Dߗ�iT�G������eO$[��!��<�z,'�ҳ�0�^ȉxy7/����7�v��b@����t-	1z
g�V@Tgu��7"��6LjKH �'�g�>�|2l�|~���]�M��#Q"�(x���n��π�F�b���%urF��9�QJE	q���*굮�8@I1y#]�t��G�$�v���LǓ����������CF-S�G�k�ǉ[��9��s�d��\�W��V����^U)�NM/�e{��/k-�UE�
��(j�8�I�D�)�yr�C�Y���{��XW��K����RZLC^əS/��4#])��3��`�S���瘒� �>7�j�o9�`�!���]!�`���w�;b��R�/-�	L�gq��*�6�\cM��1,������/�B�@��sÑ�I���^>IF��J�R{MH�J��b2p�h�Ə�M��K��\�3I+��k��YV V�S���`���B����~�H��}>�?�*t�ķJ!@V$C��:�Ø�l��y N���<�����i�c�Lc��K���X�7�����Z�Z"��kv�M[EK���
��\2� �o�璻>�j�����A�fVv����?}�#`�A桤�k�w��J5X+��Ǔk�o Lq���O���oxR$嗚&d7��1��wD��D�;+Ro�*	���{��.�I��	_巤4���NK�25��}���J�QB45Q�c�y'Wex7���ҌVZ {@YFG@�����UA�j}aГ��v�)톖ش4Nx����� _�K�oܣ���"?�ޑ2�z)�*�����i��'�$�Ҷ&�7�(Q�M�bw��JPQ�_��n�����4�o��w�e�˭�@0��eC�34�0B2&b�$F����S���B�Z����B��f�+�``�܈�*�M�c��-�$�n�0�F7P�"��t�w���cY�v�d�ϕ�1�/"2�È�&x��"o��N�DW $�|�3�d1���rL�4p�ͰF� YWh0Xk�=��y�jM��OqCd.�g�<�b\6��߆�eh�ݦ�5�I��"�:miڹ�@M+^i��T����X�9�Ө� �%�jk��i�[{�#���n'�
Hq�4q�`��6" _������;��8_���=��"�+���)2�x�pa-���Kn�)1?U�Qu����1�wm*��'�6�>k���0�(�-_,{cO�:-$k�þ�#3��I��ػ����sM���V�Ae�t���rk��z���,d6�f�I޹�ͮ]+Mm���5U@`��D�xZ�5�r�}l|�����*+���h����"G;8i��>�'O��E|�E�-��?�T���#.�G&��u���4�u���+8�_�Q��K(�i����n�X������,h��B�钖]�Mf����jQ1N,��o��R����oj�u�m�yqj$�R���'Z�̣\F)F�,T��o���i����.O���Ό_M	��!�^K��M{GQ�S�V�,ݎqP_�/LN��un�!A̅�X�+�����w���G��{%%J�0�cu�����a[BLL�Z���/���k�Ϯ�Sbۮ��C�
�� 1�K"&NX�ƕ�c��F�Q��0R�����7�^���ow�b� �Gź�_�s*�aK6��w�Ĭ4k;��:�
��9�s�^�ek��|��WMgg�+$ t��o��|0�P���;]Z��MC��s����Zz�����ϭ�w��G|8[Я�U��rƤ��q���_NS ؕ�nnm�hł׎�8����Q�ىm��F-jj:<c+hCUc7�X�|ɩ�O��BV i���U��!�,/�w���$S����P�����BL,^0�`\/}VUšg����c�np�B��#T�̀��&�I6����0V�NղFU�0��8�:�n,�͒����rGH��U����?�u�c���m1��9�􎠷����쐲� b��4��˷��h�O-��%d"yM��,�cj.sݏ��3i������G�� ����[4�g��X��Q��`,(�H$�3-�\�?�t_u����S�$Ue����7�����)q:�f�0���h�_7�#� ���*XA���|j���ľA�ܯЖn�w����+���r�LUKL�	s�ʦ��KaC$l�҈�
�yv������
��a����F_���{{Ĉ�{�ǡmg������E� l�D[z��2�8�	S�����)�Q�?s��'�wz�y؀�$��*�)	����
I��d������P6��I���>�9%4�G&Ћ2mnbEgi�g�-yC#��ȩN[($c/N��p&q��(��K� q��O�OYN�=,��g x􎇀�X�p�v�5�	p�����s{Z,S�7��k�p�@(R��e��!�}�zÊ��C�b��]s���B�lw���<�_��%�P��'��f�hQX=w ���s���^v�n��CTӥO}��d�o=Ø�kqR�������.:�D%�'��0����)���g�i����A��JU��`2��g�i%3ca�|�D��hu��kCN2��)��ї�D�����!C>:ߓ����9qv���j&ѫ�i�^�wC��
9�A����?a9�}#7l��?}�2�x�j�ð�d�ś8�G�q#����O�r����'��Od�o��i��>��q���k����%�H@+ ��,;2t�����BD����g���\���z�O�r9��F�������E Nd����-l�Fj���x4,a��)�`I�Lb���zfB�� �v��8( ����_&�!V�ҫNj��nIhL��(�> �Z0_��c(
�b�m%����j��]�֗�lDp��ˀ����m'�kY�y��i��>m�ھ�S�S��U�5�tk�r��K�)E��7�i�_�t�"���G��T�
{����v�o�^��A�X��;P����AC!Y��E훁h>"��S�4�#�՚4#3�)�h��ͼ���l.�#�=�!���A�5�%n]ͯY� �%<R�J�.��9�#;���`��=����漚�^S��=�[�B��/xp�L���2R� m-�<}|Teb%˸:W�8ݯà~X��ԧZX�	�̙0Qp(�p� F�g��m�[搌��05��&>L�����g+����۵(���޲{�*�H����_�6@���z+О&in~�$52LE�����}����|I&��E��>���^���5�Q���H��Y9ZbU�e"��}��$��k;,pS�h�(�˾�;�p��i�Op�rluaiۓ��yL6��}�`q�d��6��bH�灪��r����X�� ���[���Kd�I��{��XKd��ۓjj���+��� k'i�^	'+Io�"�޲�	����y��ȍ��\q�O���W0���Hazڮ�X�ţ���]qC�����9߻m�E����` ���X
��K�Ҧ\��z�`.g�a�z�w�&��}M~&yy�1U�II���u��pyz�7/��[֎\�jp ��"y
�#��&��hcު�\����]=�n�D�� �ݪ���et��VЛq�7<U���[m9���Ue��}�]v��#��j�|Y�� �C�[�.�����9���ï��{̻=��?s����Wc��r_?V���" m���f�Wq`rv?N��5���|q�*�Z�,g���r���j���-��d�<��E������x�!.�s��r����x���NH���"��H�Y%�+-qΖǳ�Z]#U�+�BX�`�!�(�v{,�հ��v���n|5	�l��:��O�r[7I��7�COZ����ЦΛZ��6ݺm%��D8���o*mi.M;������`��m"
Ѱ�]<t�j,q�����
çqtQ�Ls��uA��}\Ǔ�4�%8�((�?��1$��SLO�	���qO׵�Bؓ*����,jG�'SMrV����R1JJ��������WT��g@b-�wjȞ����.���S��&�,�y���~+`Sg4H�b�����*�S��0�R7��p ���d�0���5�?�a�_�bOS��[��͹;��ġ���ڇ��2b�� �fX�%_q�W��t����MG���3���0�p`,��6Vgn]!��p2�҉�#��Q��O>Rq�l)�ȧf��:$��cOo�p�S�m��C�p�O�}���wxI�hp�c�$��0�ˀ��@��k���{c����D��X��9ҩڐTUR�3 ��`��o6[ Xo�0y$�cD�����oE7a|M�����KW�*���ڞp'��&3�h�d��#P,�y`ꝼѮ��4��@�0C����I�-U� �c�j���m������s���4q�5�� �en��M:x9H.�0����N�?.�,�g����Wy�%�W;Dl����#��m��6�5ا������3
��h)�,�~��P)S��_N��rI���U��: Kt���������ȿ�������J���IL����(F�����~$'���tv��7䓽�)ɣ��K��M`��I��R��a���-`ƿ7vܪw�a&�
�o��,�����|��(/�6��SR�����V3���̇��"�����&�	u噗����Nu�ԉ��K7�-��l��#�ĆP�l�Ez���*:�RY��˄�6AZx��M���� 5)��ay���wM�#�b�Lֶ�e���9��ͷ�o뎌."�zSn�1�2"�j�<��/Fzp�}ճ���2d��C�{�	�P�a%@�����J��!���uq^8�"@��uF��Oz�(h�W 4^���~���~���<�!���F��o��<+��FC��#�0a��Lؕk2�i��{+9"y����溮U�ce޿�����MǨ���.g1��:f6���M�{1�3벯,�.o�_&������I���}�K�S����e�p�>�]}z9ه�P��{��.�Q�j:�v�)�����G�l�G�%�!7��/��[A��}�vJ����<!:[�K�ՂN�L&&A�L��O�`�D;���"�w�IY8��t�����I9M�h@2u�*��7%�Edsʓ��u�v:/��k��^�R~��P��w�Ull��C�U���ΖZq�<ò���\mt��W�Y���N=�)�@��]u������7�%{�S[PLzC��D���6_�%_W�2}��;����&l
�Ԟ��Le�K��B»A=�%�wP�	���� ��(kp��@�+��FxP]�6{ �I�z��t󒬥lJ����%���v�f.��z�o�k�P��a��%��4��*��,�i�Z�L�.l���v�S"��4�������-m��TP"�ڮ"Al=e�29�鼩�#�\��6gT)(c�]K�����NH��æ�,�[�X��,�� /�]�{}
+R�5�>���,��C�tɇ�ة���0��m� {b1�l�Ǎ�׽����U��@��,ҸB�v��Ia�""?���@iؐ��><@`n�Q�h4�a3�T�.m�c^6G���ӗ�o�}ma􎦮��aX��n���H�^A�U�۬!P��u(h��U�4*��%��`�X&kP�z���}ţ������x*i�ۥ,��6Nj��h�ed�~8���b� ��ME���3��>)vlT�z�YP�Iy�$W�>`�v�[/��� �>C
K��Ak��r��H��w�!��d����eޏ����Γsg�",�̚��5�*�{Sx��^�n�d6�u�[o��KՂ�|:@�~��z4�t�,_-���,t(͖t6��T'N��+5���,�O-%B"�����<}��vq&�H\����lLa������b�P�x�3���`��4�L��'ۣ���A�W��#8WD�$��aP�Ã����P��� ��UGj%��&�V���Jg�.����Q�3�5
3"��p�����-(���ӏ2��Db�q�36�|����ۛ��Z,5���g\�}YH�	��}�O/"R�]�S�9 K�@!G�$�v�;��75��h5ͯ=Xx����< �+�G#3X������1�~ʹ�~��}�g���erIb�V
��, 9�F�
��s'/�\K��w���̸�-y(�Z��Mr�IO!Zh�8�N? ��kK�&��Z+���ڄIT6mRC5�+qc�>�Bk�^Ӡ',]�Ͼ%��Ǿ8�廁	2c���R̕]��{�|�d>p� r�5_������3l�4��RJu�y<Kh׊se�`t�'�X"��2��vS�\�֍f��q��"X����V��Ԏ��c��aC����ŗI	<�	��XY";f��s���:)g�M�A�I-�[O��y��C��C	&��Y%�x>�33�V�jܿ.L�I�Vu�֢�+bs�>��o�e �4ّ�����u<6%8�=ޏBkc:�p`4 �}-�T:Cy@sEԺ!�Ra��"�F�m���5R���+�vԶ)[�h:��(�n^��a;(��7�vz����N�j%��� uy����#�lc47N%���c�X�ڎ#�


�v�.�a��a��B�Gz���Ғ�B�\�{����4�����"kY�=x�O�(��ۙ�2qǚ�=��G\�j�y�,�",�v��<V�O�^�c��|� ��+gt��w��DS`�?�����h X�j�<�XE`w�?���-��y�h8�K�>z��1'�\�M��3D�\g�����
�t��^^<f^�Nh��������>����C �ທ��#��-�`�=5�b�zK��Z)�o�EL���F�U`�w��r�J��65���RH����r�	>\�O4���Y堓I>L2L�}���4���<����2�}���8����(��%u�4�"3��ӥ�HPۛ���ŌR���v�k~>�,l������5�)����4L}���PBH^��d7������$�9�OhJ��/��r������6B|�O�"ѱ�읐|8�n�uG��/6�i8l )U6�@�s�E�8��iP��b�Ʃ2m8����7�>�Z�v�a�U%eL����J�JX{`��s��wM������a��$���ϭ��s}�!4�(}���¨E�����?OU󳭥Փ�,�;�e��*v�[�xd�z��U������{�q�=�`�5�K���Ƕy���k��!Q����x���~~<qҬ�fq�뱵W�t���܅u���Q1���������e��lRc�)�u�Q�Z��r���D=&K^�;�z����1�x��L4ؘx.���CK|o�m�	���./�r�Y�X�c&�	!�>$��ģn՚ogZ8����c�
��b���@Ni�(��W8�90ӑ��@�3��sF'k�s��m]̓�sY�:D�Aǵ=|y�����e[�v.�����aff:�dx��ٙ&"ȏ������.�mp�d���������m�x�C:Sb�@X,dx#��-�%I=��r�T&*���s8�����d�y�e�������Կn��:�Q����Nr�Cs�?ǹ|�ZZ��~��(����oɎAI�cJ��8:�(�;��L�-Wޏƿ�2�#f0�4n�@���l�M�!���f)>�~뉘����ܝ$J9%�����.?���dz,j8o�y����hlJ3�+�4'm�27�A�0���	ٱ9=ykb�5�&��ه�?�����	���O ��}�䗔���%g}z�.z(�RT"&l ��G��p�	o(K1��ߨ�A���̑>3!Kly�4H���{�_��$�6�z�e
���,�������.b���vZ���`"f��sX ��)��������Q����N��B��ftb@�Ct�t8�R+������e�ow=�g�C�.��"�
��r}�`%�G=�8�᳐ݴB=�����njU3�>]d�̧�>�^������9e��\k@4��3*\En�`Ŷ\�w{� >`���z7�;>�n����:��W�!;{����h�>M2����vN�;Q��l9���?'?ޔ����a�^@����&G���j���Y!4��&\��R8�^�HVR��)���SS�Ro
\���G����G{���@x!��(����ڠapZ;cX̶ٚ~�	������B��BC���NxA�at��O�e��c�4�l�sGG�c�[���n�o+���D_�JC}��|����Y��LJ5�C-��H���-�	9�gr����ޣ�l���/©E���!���oP��fNz�OW�q�˖zΛ��)�!���RW1J ��>��Cc"��iS\s���☗�w@�v�g��8ll��N�'}z*/�J���Z\�j�/窒�\�Kһ#��ɛ$�r�(�53��W����T}�Ű-P5��Yc�;�R�k1���)�ˌ/�N��5�	Y�T�UF��W���A� [PWT�NP�	,�����F�ips�l�N�U���q V��_����b���e��D�K��A�R��|op�\؃�����{ק	�/0w��ո��U�,�z��4��g8�Oz�3��X5AQ�=��{�(UYR�_�v��n����G�hD�Fu�7��V4�KK)���yF�)	�XK��҂�V_��B�H
�$��G�-o�������n���$M55���U�Q���ݔ�Nɞ�7�삯B eD�\�X��O����9���D)8n[{G��P��k���Ãf�W��GM�48;~��o�j.lǡ=WK�J%+vh-�IO�3��H%D�w)\jlQ;s��ݛ>�MO�&c�o�Խu+�b�>6�([̼��4L��Fv�̯�K4��,J�䘻�&2K�_d��u ���!�Ĉ[������.�0�ց�Ъ앗��,�k�e��7�O;��=m���c嚽j�'���잋��d�p�K���	�9�f�G�_�'�祉�D��p��H��P������K����@9q��F���{�t�xFC�z���r����J��W,L��q}�OD����k���u�n���}�hU����)���
��M���Q�1I�1 �0غB\�|  ���D�����2_����Ĺ�C�$ж�779��a�2&y�~���Pf���
�ͬ"�dyG��A`���3B�&;!ˡ����Kz��$,x��ju�n�d�F<�l%�p��?�v~=ߌ��<�iyӱ�	j1vˇظu4��(q#5���-Á RH����El����A��7q
İ�_��
D^��v���4O�=��Z�!*H�F<%����lC����+r��F��~P�R1��s3�mA�')(��MeϾ=��_�ȳŤ|�Ǻ{j~逌s3(VƟ������-KC	��@'��V���P� ��A���Y=��h%>�Azx~=o]"��?	���r�6a^j7�`�C	�ƝM���1L*n\f�'k��k��R	�̽]0
��Ƹ��u�i֤Fr�)����r�:��~}��,�6�s���6�a�D*!Li�L�L@XU�CR�:��������?�^���آ�Ys�Y�8��sԩXW0� ^�:��P�+Pf'�T����Ñ����
���_�%F�2M�B��,`�x�S�;�`"?�%#�Fn��I�nO������]D �yd�kſ5����;o;��Ō��n��� �P����l�yR��M����S�F��>���G�l8PY��ʾ�u/�����g�-�`u�Ph�|Dx]��<�=��9�}����f����M��_�9���$@leqRSy��<�0�^-@������	{�~�������
���ٿX6�q��q�|��Lh��/��*��T��a�H%bn�*u!�T`�/@� �q�\(�#��Dr��U�!b�4�<A�'ؒ�H}���a^ɍ���ySc��{�΍�=��W�?�`���1ʴ�h��my�0 �S5�ĕQ�F&��..�0{�F�?��}�F����D�3:j'>��Z|����aJ_�j���o`�������eΚ3rCr��U�	&L�`�P�I�,2'Ԯ��M����¯.�(�R���1�z,O)���*-!aڽ�$��K!!��C�+�Cq$��Ĝh�&2�~kfZw�]���kC�3��� o\��.FD�}b�%* ]��&�$�����T4�qFs����+��h<��){�E�����I~<P�[�����0��u}�4����1�Z����%��l+�W�A������^���E@�~�l��G{��$��8�T��2S��"ګ��x@W���C�����vd2� 9�t��g`�kӂCk��f!�a~d���uMY�i�1b�*�~��Mq���q�,P�=�4�q����۴{��T�N`�1n����y<��g������A�̈́��l�xv�*��0�Hp 4���	����iQ��V�����%�\���J�����a<6��
�E��SZ)���z��>M�A%_����I��+6u�'�m��2*̣П�e!5Ç�sii�ܞ9J������IQ�]wȁ�qy��h](h��,����c��@i� ��9�2"Xut�/E��X��|��|240�_�R� ��o�}�9JMH��ϸE>B��m�!���2��d8���/Y��p���*�� }A�fq����c]��3�(ʃ�aV\]oQ@Ʌ�N�#�M_<ڨ)]&�&�ՒI)^�e�Q& ��sOq�D~U�Ūc7	�F>���uA�vK_I��'�o�>J��������1��!��iU���$[�ph"vַ\l���$c�`oZ�E�ۦ�<p��|�77���`niA!(��/���o�ک%"����-cNv�u��l�EDP��d�q������="h��g�M��7�z��p%"X�� ��Z�T����w�\Fo�it�/�x��&�p��%��],����B�g�I��:�����2����}cTC��c���I�qc���Ó��|�����@�E�L9�f�'��jA��o����nR��ƪ,	'����O>}V*�vU��}�ɽx���P#p1y�cdJ/W��~`�p�
;�X�Y���e�b:EP�O���%��|�?�#��S���_��́��5�֛&�ug���T!g'�[�"�5*i5�'��g�C�lk�����B}LQL��[g]�ݞ8:߿0��
�걛����[���i��,�ӳ�gА caoښ����/3%�?�^/��q�M�� I� j��L����PI?�y\s��U>��p(�Gy���Q�,v�X]�bJ��ZVw�sP��� X�4�(��L���eP��#S������m�L��"�e�;(��%���X�V-.���c�#�nl�I���ㅅ0�ni����F���U�r)�u��xIH Rn��+*�#G`��R�Գ.����$�[Ʒ���@��������y��/��r'��^�]v�'ɗ��0C���(�ܡ�#�
�i�^�mZ��d`�1��_�m�g�4*���J#�����7�$�K�[�U��Q�-׭B�:���:T�
�������+GA�(�	�@{��|Io��"��f��9�Fg`��5ff����v�~��������f�'2}3V�s� ���Ay�`sM������B�.��䦳��
˱΀���e]P��('b�/W E�=��})�����"��6��/ț�V1)�,{���c��ܑ�B0d��u�:�H$�����t�B���/�����Й��v.�7��n�G9��\���[�<kQ���F�
���Uj(��X�[�@�7���,�azf��ci#O¬J������;b#=�x
N� ����;�3!� ~�^���#�oe h��C[�ŭ����} є�o�:�*NL�g؂�m6"*,��/�	5���i���ߚ�,��o�U����t��G��bٟ����$����5Y|���Ԧ��NA�;�Ӗv҆��^����v��]<�q#��������d��Z�O��-��jƜGn@J��ٝ��bٚh��,�
���X�B������\$84e�Y#�"���YG�-�|��� ?�/�0h�a�	�6iK�� �=�fW\���{uֱj}(41̉�+��-�<o�������/Ґ�2i#Y�^��36с��	P�7Q����c9�p��Ry5�kF� �S�b1j)eG�뱟k�����b�W���(�9���`%Mq{�~i�,��o�KLZ(�!��2�W0O��NF�>��J�T�&���2[$%�r�:��?���b������^&V�󑦧E���D�I����l�g/{�$�^v;f�b�8B�=��p��� ¶���N�����7�>�`��
:lu�Hb2J�A�J��;� ���
Q���Kn$F��Y��ew�պjX�+p}�.:���r����t#��
N�j�s8Z撻��VD�b��V2���u����4�-QeǶ�ًD��^E�IG��Jp�{6~��Ih���D�6&�.ɉ��y�z��(�N�Q�
��yf��BB
$��29b��&z�&l'noϗLT�Mm�G׌��֋.��l�u��M���Rͨ 9_wȁǽ��h*A��z˲`[�$'Y��Ь2g�[��T��l����oϺ >nZ�JL��E���I��){�I�@�ǕUagI<�K��%�)S���Yf�Zns����f;*�Ɓ-,��Vr������]��8)	�x�,�k'��ND�4�9È�0�@�>�w	59"I&��r������]������h�Ɣ��o�^� ��-'_�xVqx�DEc�E�C�:�u�͂�}��ﳴ�'n���8��ײ�� ��3y�4��&��x�@�蟾P��<�������r<I}Ɨ��H���KcY��֮Y�k��Q�Yݔ�/0|����K���/r]I8�˔u^�el�q�Տ0/?U��[�����z�j=��5�:�de�؅K�ܓ�*B�q��2YRs-^U�`	f��
��r�(`�(�%4���?*�U��xga�|2}U][���T�Gg���p"|'��f�ZL�_HvE����w�s@a�_an����L�z�W�|��U����=�L8B��Yh��#'�ҭ9k������*��6�w��B���L��F�!�-]dt��f������	HE��7��Tە.Yd�D��F��^fP�[xݭ�Xn���`w����#~ n}%^���`K �ST��i1)�-�(�g�8��?��jy�`�5���ɬQ͌V�f��!�\�,w��a���P3ґG������>��[m &�Q���T�kc>+�G��`�S^��S��2k��)���.�����}���,�����vڥ6�]h�������=`+��7�ʟ]�<�"}�;�n�ʙ�Ĉ"ʴY�~.3/7���ބ��(ݦz��H�?�v���+�*zӝܰ�=�D_�y:��x�8j,^_<;rÅ�i�f�~7[e��Ԅ��w�w$J^!�@;�h�xv��Ԅ]�˚�I�P���Qu>�Ѣ�B�CC$�p��������zo�;N�)�Ni3�U4��$�:�.��6'
J�^T_�2Ϫ�rHz��~�+r���2���	��߽�5�	R%C�e�T�R&�`�YR3Z���A^���9�i�Roԭw�X(�8�_�+�����h�!?9+�s[�2Dj$90eۓPݨ�����䥲T�����`N�VRP��=�Ñp��\H|Z0�߄lo���e�ff_�JoE>�U����Ð�H���T�(c��O��K<"7R��F�ס��[R��A�������m�P<�M��Q��ظq���|1>�Sp#��ǡ�b��/�|~��]�0����mK�и��I�T���s��n^7��L��WU=-��֐\%��>*\klX��H���o]̈'9QL�ڞ!T�\-�pu��y_,'�E��7�]�EHC��D���"�ٍ�h�w���k6�k=J�Ǟ�4E����1;ž�q�	��fL^ƭ~�(0����D �Zf;��s���BlQ!1fyƜn}ٰóLa ��2�j��i��q�c
��o�t^>6�l� �m<�<l8��txҵJ��
�W�;�
p�x��� �È�����#Mp�K�����Q�Ϻ��Rƃ�pc��qs�R�䞉��Tl�la\er�k/�������
-d(�0�y�Իa��ϭ�j�/;����A�W�w��m�F^l�U��;�a���:O}�R~�|-n��WVñ�yU	Ѥ�hҮ��Q�D�����<�0$2������&��;X����KX�m�=�y[��
^�cV"l��}<�Kq
�ѝ��v��4�
��v���h�N,��>�/^�O9��ϛ\�Tr���6֡�9�s!�}	9x�E#�H���0���+�]+΃�p׏��4#�.�E��u� �y����i�dV�C6.��c�ph�~�H�p����K��=��<ɜ^�]��a76��浀���H�#I$���Y<-z�g��4��I��@Gp�"t���
?�QKӔ��Ϥ����/���2ZLR KLt�ϥ�O��l�v#�Ƣ�a�/g�S�O}a��bd#�9��9��EAP�\�]�6�%��ĭ%�wټ����-5�E�Q��[R�ώL�Ee�"����
v�I�"	�p�
^�\gq�w|!}�dt���U��&M�᝴O�{�<�}��&��ӷN�#ד+hOkK��uQg�7��Tl�9Y�O�fқcݒ(H:��-��Œ�]���1���M��F�@}�vNla*b0�|��p�X�oP:A��I1H��v�ө?_�ő,�R�H�@_��~X�9n���eTۖ��q�X=�F��:|��<�U^9���/~P�A��-p�������v�&귊;ٱkh.Y��E#�X+�2J���󸺽O�	��/yu��ޣጊ�v��]~��5��u�?;w1';���_��}I�-sk����&�=8���hǥ���+�:��O��,�7})����`g�p�4���Xn|)��3�`�k��j��Z�#C� NU�՞��$�K�ʞ]1���3����L0�Bc����Ȓ��7��Ҁ&�ظ��{=ܶ�P�s|W?��@�x��c�[�!	-���쥯�l0r�]ݝ������s(.���+H���	�
����?3������|����(�Aނ2Ӌx�2a���!e�'�7˒�ț�ǉg�J\�oi�GƏ�\��H�D �y�"sb��������Lʐ�i���)�x�]�`uXC]3껔+��
�	����3`)�!"a��o4!/�	<]b�������{�<�Uj�����}�^�>j]�ܝ.�$l6����}rZ�:�t#p���,"Ɍ��>E����X��Q i���O���S�=�>v$���/��Y��}����`$�뫊I�1s9>�W�S���گe�P~k���zY��;0q����6S�U���45W��i
v��'Rެ'�����h��I#�.�b+��C�=4n'�����:;��L���lV�����|���x>���k ��R���&�Ar�^��t��)��|�W����5:���أ�ƥU�H����А?2f��@i̱�/���M~WYxS�����R�P�PӶuze��9�u�}���,�B���1���(�L���ۺ�n_�c�1L�Tn��w�FZ�G��#���8�P�԰C^!jf�ڥ��kkL�z?�M �8�L��iTcRs�!�|%�ΒϽ8�]�Z-~0����$���xZ��ndD<�'�G{|/�\6������C?Ea�`�"��� ���P�rI��f9�ե���[IA�=��1�/[E5�je*�����Gd�����_ᱮ��;3;�Gc7������1�m��Bh�p�9��VaJ�+�%*�a揼�t���'����lF�葋�f5:�C�nrg~�_�`aM�G�=$Z��nf�$�?�3Z]uI���	V�����KE���\^�c�IQ�]5ǾB��7�C�(��lw�9+��M���uXVbL3^X�C�=��Q��^�ܬ��� ���q��h��M�zK��U;N&u.���]E,�v�J�%��Y��'�"3����=��7;��GԫR1����?g�#>+9�kz޹J��>���a�r�t�]��%y3VY�	���/0���u{��D�mؙ�lYYoT�þǹ)�{������=.�'q��.�Rf7���.��2�1�U�Kg�º�Vi=���y�#:�����M4��
&$H��{��tL�wLQ��Ty��Ƞ��� 1@�@�q�*L�aH2P���V�}ǕU+�}S3[�ٝИ�� ��f�����4�zĳm�2)=>7��P��^~J��j���<p�����c��5$����[��~�"��TD�oi�Z�,�ވ��.��$�j�:��%�a�Ȅ��8�0sG�0/��b�

��F����U�]��(|�'��V���w��� v9��"�p¼zo�EL���~ TT����2r����s5S`҉S�<���@����6�e�`�-�Mm,��f<V:�Z��y������1;��#�퉅�q ;�s�΍�,]Fߜ�I�_;�r�e�4���M�e�"�حL��8L��C\/���=(�3�x`����uN⃃)}�!�3R��Y�'�b��z�ƬfV�!<4�4��QhX�O�+�/�g_���ui���f4��@$�g�(�1A�a�.�L9�C�A�F	`�*��3l%/�A�P���BS�~���_�3'�'��ҮcV6���I��2�!����4e٨S��(�9��wz~�{N`L��]�
&�2x��ӕ�S3e1
i?��?RA��:n���m�k���p=�@ȱD���,���.y��0j�q��m����|�T�T���<_�-=��`��n�;�Wn����	��>ˑ�o�����]p�D��,�^9f�G��~t�Eh�3�h�CK�Dڒ�9p{�?�ڄ�b}k�f�s1����]�}�6�������o���	~��d�(tGH�fti����ު��S��q�V*m� U|
��}�/�I�y�P}P��U�x��=_M�R�H`��o���2G�W8��?|a�{�%����Jk���n.�ղ`���vܰ�����s�+�S�$v՛��`ge�pa��t}�0��F")r0�_�/&o�>ۄ>^�4����y���!�7ě��4�o�õ�����f,Թ�]��J?0ʛ�mKA�n�b�m!�G���*��I�$�8(���<Γ2�ji�y�l���G%r� �����S��������+�p2yv'T<��>�*�0�	��?�P��$I�̔N�ᬒ,�R�^E` 1���B��ܥ��jT����j������g��O �� #��Ō+������h�l��Ԁ�,=Ra����lx��Ml.�/�@�Qj�#�L��?�(�tC���?�����azRQg\2|ܠ��XC���~��@��˜�.��r'�X}S�_�ED��Ư�]	#�a��"��2��;��Ԫ[C�U+��L�g̏�nox�qY��	�	��8a�x9��o���-7���<6֊t|�ӤEo���O���pI��E��>�G
� G�f�����2G��A���1t.�"p�q�o�������ji�s�:g��+`�)䱶�P��_���!F���rJM���MX_�&3������)���J;6����ׇ�G{���Ǉ��;˅jjMr�:Ä>��5v��$m=� ����;���O����>V��+OW���ɛ�[��`fH�+�a���&Gjr/Zr�kM�Z8~p�ji\��x��ap`��־E����/��%u�H�})�ıF�ylbdR�I)��܀�54�O08��r�8O����J�hgB(!?�U,��1Ȥ��n�UW�fu1�����I1:�J!�����ΖwG���r��=���� =}o�ʈ����Q^J������Y` W��=-hO��O=%�9��j!u`L��2�s|�XO�6�^u7��`zB�E��YSh,#&��r�7�	��I��(����=;*|�Ӻ[�Ӕ�cY�h�d4��9�Gf A� +�/!�^� ���w��P�sf�P|Ҧ�Kdֿi�;Lg`�a!�(�3��]�8~�Z���xa^*�T��E2������Ic�a#x���A��2@��co*~�V�amy]M@��X}�/��X#N�j�����e�+5*x�Qp�6�E�^=Pb��{SH�Þ��
;Wa+>�\�ȷ-]ib`�X��C�V �]�4�E&�3���Os�
��A�����d:[�?��i��䈦v��m�<�����Sz���ӑN�X�5��ǔ���S���O��f&��`NX��wk���ۮ�}����F��@�%�H��9��N�wrm��0����J���nM}���P�1����4Lm�f<��]V|��������}%��9F��tR�mU{�IV��1�Q����n��N�C��%A�F
?J�j�tC&��6U2E6�	�?�
E�M�k���w%� ;�oFp\��A9��YW:U�Yg<؅���,J�����s������fm\mV�Pml\��Г��&���Kވǒo/�����ajĈ�(嶇?�ʊk<6����Be�{��6=L���Cl��4��c��բ����^FK��6�\���B���pqx��;�7��=pړ�Ͽɫ�������'*M��95q���	>.W�f�I�q+|"7��^�[���V�-q�Mѽr΅��g�K
/�NW���Tȥ�~��B���K2�e���&��>c+���Y��U��ѭ"4LAG�A�Q��ͥ�a��~�3EstQ,�*s;�B��z���w���<*g���S�/u#/|ĵm^�{�o:_K:P�W�Q�L��I�ꗸ�8|w�i�b�ϸ�$��LM&[o�YJ��+�"8(�B̿�ro��ؓS��WO�q�K��Lt8�����(W��xE$<�[�k�C�u��z�վ�64x�V�${ SM�7��i)�r��0�=�z?���13T�+8P�J����13*�߀���g���`KEj�xѝ�[,��4G4Wm�>��1�-:T����P0Ƅ
=�|>H�n�H�9��X�/���N�$��x:�A������"�#���3���j�h1G
{56��dlǜ-5�>Bo"F��2E����I�*.��c&�7����"���?��c{��B�����N��,*q���Z�v���/�r�ZJq�"�/�30x
"�r��9��6]�5�t���s+�G��浼���V$��F��0�?>s���)��"�sm� �5���6�݌&F���}�iК�M�����?���j���;X�P[,Wu��v��sg
�s�\���}�7����X��إ8��C-K����]�1��E6��`E����K$u�u�Q��A�"�|���k9և��ݍk� ���̪h�H+�
FS{�8�T��
p`'�V��I�%@!��!�^u��%뷧%F�{�B�G��z�0]V]` ���b�F�L�m��Gh����.r{��(2H$�I�p�^��:����J�SY�ԕ�J&� z��R�;�	�����GK���D@P�� ����
���2"�4�]Q�YD�\�&mrc"[�������2M,
�&���-�m��k��
Fe�w�4��|Y�?b�w�p���Ǭ��R�ܐ.԰P�ּ���Nm����V ���\�1���)� �YO�A=�$P��T(��*��o�
�ʰ�h�L�{o���/a.��vJbR�6����	1�/��d���cq����&�|&P��9,�� �p4
��b^���څ4m8�~��
F�0�̃�)fW�>xp,�x0�#��Iϑ!��3���(�Wc_��S1�T�G��q�������u3�	�'�p�iA��n�����Ϲ�'�ěgAd7�id�$�L��P�!����i�2�%�'�W��s�F�4�G���h�X�bZ`Zf��W�u�:/X���N`�}֪��R�7��������t���Q���%���&��v��l�|)�r�8�i[�3Y஫��� Y��b���[�,��2Z2��nw4��l�1��JM�SQ^����>�<Vg�[y�I���i1��s >``x�k�_� y��\���i{��&}��&m��x: ل���W"w���ԗ]��dv��)KZ+�MN�/i3�s![�z���9K7+���⨬�����;�����@d�D��M��?q<��K-=ο�e�k3)b7/2^�^=�|9�L6!��Ӯ�,�G#�+d��AsD�ɷclr�O��?X���M�����t �J5�}�\w����|�W����[D�+|G\�t�@vX���������ۆ������4z	�!��F)q�+ً�pfm;�ٶp�L3y��`�����;�ɽ���O������X�Y�Ц�i�!���.��^!�݁~�ۨb#�)��'4,N5�)�X�ƹ��ht�R���]�	��'��-vs��>zų�?��A�������wL��i�{�@���J�J�aW��.�^e�~N��<���s���.g��4�^C[b�ܢE�Z<�@��6��t��s^������'����%�(�ީ�Z㿇������O�O���2N�91�0���x���k�5�s��=P�4��M����� )	�r�t顋�7ב[|�2$hp|-v҉Ǎ�9�X)ns@��N_���'�	j"��қlۘ���� �SL��D�����t�̯wۓ�����ƭ��
<Ye��7���-`̡yD��[�2%s�R�Z��ϳg��K��V�v,y=n�U���yq0R���� ���8�`� �5ޝA��a��Q1 �d���F?�?>n8���3�d���)�I&��<��>T�0�=) `8��=��oH�B��܌�8�g6���"�(�V�T����/ݽ7%Xy��۩��~�Y/;��<� ��]�>�N��E�9�&�x2���i�UpJ4�F�����G�*/Sf��dM�1F���yW����<�搅[�y�-/C�1����p��]nZE��xj��侯�����Ϻ ��ɫP1���(�jJ���`4�*�F�_����7�X���.�,�2��x�<��L�T��+�m�����U�Ge�N�y:���l�w��&'��WT�:�*6@���6�8ep�Q;620u\�*�S@'�_�	CAf��0�]hK��ho�m������WBo��h���O+�LAy��P�13,+�K��%�.�S����L�$��Y �dRf�d�U �����"&��O��	R�â�tH����£<�5����7sg���p��<��4y�3�">D����I�e�~��?D;y_������&�{���P6�,P;�6����&5L� �ƀ�ݥ�aN��$�v#C�90־|3�0�袶:!-���XP�v�L���<�u����<v�KM�� ,7��4_��ie/��Q��A��bz5���XS�O8ߕ�(i<�N�*�
i�z�T��(��AiJP���h��V�����s4NV{�u�������]p���_Ζ"u�LB�!��J+39�0]$[t���3���!A(���1���\�g���P��8��i���2�^	R��q$]����R����*8��U���-팏ӣ�h�%�j9Eզ`8�:�Z�,}�2}`h`����ݰ'<�������Z%#��b��%��D�,�'�,���O�»B�Z�;��Ϯ,~߱�~�E��M�@�.�wz�FRuJ�9��j�;yÔ!&l|G<�>۬��1ϟM���F+$Ɋu}.��F��os5��$�u҅F�uɳ�*�{��f�ٿc�Z�D��p쀁wa��I|�a��Qv�ӳ��&6"Gp��?�@p܎��s3��@��,���A�*�ٚc2g6ʫ.`�ٵ��9�4e�y������͍���M�����\!��U�#���#�B�}zk<�+j.ԡ�1o�o��8����-��5�k��ʀ#�_s��gd��և;�`�z�f��/��D��G�r��h��ў�d�@��5���+x$V�M�ߗFJy�â,������cFp��Ss�{m��4���[��b�B#w��/}�=���}HR:#�S��#�O�S�Q�s�'5����B�8$�p̆J��=��&A��?�K����Pm�h!.V�;,�-/�� >POF8��4��s��
�����������j�80�8�п}�����G7����X�Y��ULA�)�A�{�&�|��ʧ��`q��J���R�L!cy�\��W_+��_�,d0����,�����Z�vkЖ��� u��$���)����Z�N��1gK�g�j�C�b�<M�q���Z~g�y�w\+��;���E执����4�iaq|3���H��
�F�/A�}iI?���m��=E H��N�읿˹I�O�zRi���C{�A��2�w?ֿ����ǹ@?or�MٿHk��G�_��6A�j͠�Pz�v�AY.n(��O+�`$<Q�^��f4~�0��pk��}M1⺺�f��p#�N9�����=��HԬw.<�����y ��.�Ԭ�Ej\齶F��=�V2˼l���;�\{{Sy�Wr*4� -�4 �rh!*�M�/7F��j6�58�������꩎��^�BÈՆ�3!�*���K�s���N�NϚ��q�-X����t�l�eO�ň�N��y����pfa�
=�Y[m�S�E���AO�`�2TN!��`���6���<X�@���%<���������`�N֊�Ut��mD�F�/o1�pH�x����ߙ��t���d�����j�����J�6��<�{K+4�ǀ����r����e$������h���\3S�$���>.ܵsb�:�b���|t>������y�������Z�n��k&UM;�؂�/�i�����ߨ9�%�*LQ0�/�_���ߧ��jՖ�܋�tp��gcӴp�H�4]�[�`��ZM����:WM�k4ri/MWPgV$�=bp=v�Y��ۑ�9;S�l�����"&�z�j	D͵��:���*�Fq��b���U��3&Q=Ŵr�5�JN=@wz��?�ֶ7� �0�"~ۦgo�hή;gb�ñc6��h���P��p[S���]U�tY����x��ٱ����zh!�P��c��ϡ~�(ܼ����a�hg�+˲]�-6�_�D8�3�{�k^V�1�v6Wcs���7�_��D:�J^��r�0�1��ץ�<�K�)sJ�� �%� �L���r�O5+	�"�}[B�.o�^W,�ӟS:�)b����F�@_���Ң�6~�J��Y�A!vҭ����U��4hp��cV��Ϗqt�Y�����]u6S�T��S3����2u��~
�?������`��[�p��g��C�
k}�Ӎ��͸2bS2belh�������sƧ���������+e՚ՙ�f���$�Ea�C�"b�~,&�<jc�6�2�kK"��l�8�� *Y��v�N���\�W6��c{�W�	C�o����7_���'L{r`�mL�(뗊�9���w}G���ߩ�:���@j�Y�;��@�[������aP��DD��\5N-���TRqOق�G��%�Ȅ|Է���`�Zw	m�S�����K,C1Z������y��uH�8w�Ӵ��c�F����FfNx�)��W����H�0u=ğ���\_y�b��Us<_�cF�`��I��#������8\��)p��;��G�5��7�K8��-9���)��Q�E|n�e�z�PsX��RAM˰�J�
�u�.�$eU��,7'|/x�{����N�i׿x1P��aGC��� "ğ�>�#������������
�R�L5�u�D��<>ZF�ٛoa��v���qhك���ɧ$g��w+����r��U�H�(h�t[eYu��s�jV@S$�����1�=�[������Z�z�����g�1lGCW����u�$��$g��M14|��׌���ۣ��*��fvj�������yߗ���+��3)��/��!`]�.ǎ�A�
q��b�l����0GoG�5� ��.\������e�75����s;[���zI$�M����&{M(1Nl�ɻw��� ���D���*��VT���xv���.��s�].=�Kob"���=j�!����n��8wNձ"CU�-s�L��ƤY{�,���{#%5]�Cu4>P�@46[��-]�)�Ǝ����P���h��u��ZŨ0q>�f��n�j>��V��x��W~�byL��u��Ыӂ�QƗ��7{~���1�VV��'�MS]��m����`(���E1~q��#ܠ��.���r�i��u[A�n�3!"t,f(IWhUb�\90�4�-� _�*B4�9��[��B��(~��SĞ�d9���T�	*�Z6�`r9�Z�Yq��ʏ�QXAm�p��װk� z���]��� ����`�������=Ԣ�/�!���t �+1���Q=Q���%lگ�W,��F]_�Y�}m�_�^���l<?p����##Gʙܧ9�#��3N�BG��Ak�C�f�{
���z��u#����$�o���d�j:z3��9[�����j���ח�s�e5оp|(�k(��^��m@�Y�:��c���ݒ� z@��@D�aj�Z^+��$h�I�u��.�)���'��-.*C��­������=�#YlH�Y�?C@#&��;�P]a&J;���,�Q�E�<T&s�L��8X���|%AB�;�홐�ƅ�툷ي����%�FSo�<��)��~ԃ�!R���ָ 9�$n�!�2�Vf�L�N�������"��� 8�����=�(Jo�:8�iɍ�c>Znd4\��yV���w��R,vp�P�v����.�ۃ7�d8A7Ѻ��A�q���r������\t��&\���KZ%���X��	����h߮�G���2#'��՞G��
s��D�Ν=�@�p4mrĆ4J2��ù�3��~�;N>F��\���$/ݛcu�3�s���;PAJ\���
���Ojgn90!l��F�<��}Wk�<aQ�A{!(t���H�cnsu�@Jn/)�eR�����:�tZ��]�F�ڏJ���<��*.��mq���S�XɈ|�w�O�2����e'b��~�p �E�T�,0s����r�1��%�^ey�W9��uᷥ�cW��r����W��S��?F?��Q��X*�(!}��wc+�O��ߌ�:JU F�FE]� Hʩqׄ��B��X �H�F�i��5��$�I�O��M\S�j�Ny���ZDtZVf�U��=3��� �T�;�{H��I�E��f��L�|g� ���
���H&�py|�!ub��u���N�zė��,��l�:��s�����#�泗lb�=���f8N�����F�g��
�c��5�;�ڗ}B��lX�wG�#pCl����Eɯ���-k���,�կ�� u�Hr,%PP�׏8�/Es"�;�5�f-���\F@R������-��+��Nt���ǣó����w`%W�a��I�R���*-�N}�*�Q���+��"}� u�c"�������>�*F���z����@��'����c4t��ɹ��W:g�7���;��STje�KH#8B�6�᜜(#�ӜN��bs?�&0r��Ba#�MonZm��j��}:�&��H��k*<����>��`�e@D5���sR������N�ٚ�=@�w������K�-P�y���!��^�!�J�!Y
%^�[r~�.yӮiF�|�>paNAД�
$Aak}�e��;g������	� �cU��Y�7�-�5�!��i�r�. ��(���^�k��$��w]|�Ƃ�}2��m�dj�et��)���}��m��5RȖ*z��	�a�(���X��A����y<i)�� H�vnof��	f�A�KX�a�"c�4�q�AǍY���!`NhK�SR���3s����C��l##��.���=���K$"�t=���C��8;�"l�IO彷��a&q����O.��Dc��'r��=Π�9��Kߊ��N`�I��V~V*�p䩇�.�;�>6VZ����}����R���9����(�g0����v!�-LI��O
����G��0���-���ծ��X����!�b���hFQ����RM��LF�e����٣ ��ʢ�����\x���I�I���v_���#�'g��r��q���D��0���l8�����J��މO�?�e��>�b0�cy���5G+�S�o��3u6��]��Nw������ ��#�YG@��KQn�	Ӆ����|N�@���3YsQ�5`C���z��ۖy,�*�2�"��\7�*�;Hl���`CA$u���RǎkwY1q�Ν�h���Bd�P�hVw��B��J��_wV� ���Èg &Fqq��2�����3�Q*+��jș5��-9�^�.2�s��p��P���?Qfa��������V.�7&W�R������*T�ǔ��`n\��S��C�N�f�Ov:��^.�	����]�Q���E�B�W_z\��#���[�+����[28�L�;p��)ye�-]��@��q>�IS����|�Jy^�`�� J�IImR��ѭ���2�+�TW|������@"�ͩz�J+X�ert�MBr�V����f��s?0�%��uf��[������Cȷf(�J��͛qq��3e�_���v�aTVcS!���-Qw;�z�d-�E�fu����l������Q_�e���}´�blFcA���P�-����r4;r�e�I��߫�����5�G�>U�\n)�L�|��d���}�{Jv	��;c<*@�rF��t3}�;���3�DjTOщ�����h:��yRWn��R�g\���+T�������z�����JuU��E����V^�V�6��m�/}�zu��К���2W��@8��p�`2��W���Qڄ _��VQ�����Ǖ^�+|����@C�lo�7�9��Q���?~�n��n#����4Im�9��AmX"�W�4�[���0g�<s��~l��g��8�.�;O�5�T���&2��]��`�J�w��i �k�\-��L-Qx�	�d�i˱�����I�������쁐g"*��'^�7v�������50�'�"��2�)�9T)��n9�ڇ���5A%�D����u:�^i���Q��|E^O߉g[��! �齑.�GKL�H�`�<�14k3,{y��w�UH����W�����+��;�vVw���:���R9>8��;�"�"<.����/��F���=�d�P ���g1�
�ߞ�N���a��"�yU���><d�g�҂nl�%��8s|��46��Q]��@�jH�U�DZ%����4��'�6-�qm����mw�M�Yk�����]&�#���R�Ęy¸�N�\�U4{۞���Wu��oȗ�� 0_�/2��oU2��&
1�ڔ�j`���z�o٘n&�����1Xo6�p� ǀi�j�����zT��j��A��o"��F�`IN5<'<i6�	�M��kB)���������@͏SP�����xA��ӌ\��n�DY�9���f-�@\b�cnXA�y������m�2.�;��C���zTڲ8.��r�&�\[1!C���:��b^"���^�)�W�J}prS��hp��z���z���+('�@#2ݺ��g'�5��F*�e���Z:�O����~�j��A�7�<Q�FX���3u��?��V͸���~���|v�x����%M͞΀�zY3����H��/��v��<Ln�����T�G8O�S�uo,C�Z�8*�������O�r.�����/��P�r����_�\�G^'��8��B@���*~.";�a�`� >�$)��h3 �2�)�In�H�H��1&���U�xׂCm��ѻ��0���~��}P)t����pn��MGC���\��MIl] ;��
mӒ���VHT�W�W�_�w �T6Ц[7�w�@�~w�OB����b����F,\��Na.J�� D�6�<�(�����$9�蕿
��֝�#���p�ꙧ���?@�VWr�A�ͿT8�~$���}�0��n��t�NM�(f>���_w�T�)iC�z�9�'�X7���)N��U)�-�L����l��S㏬�[?M�S����O��W�ީK:I���~�Z��NM .ؠB�0C��/"f����X�
���b5N�#��70�Ȯ�Ҕ��ty�bon"B̰��@�M��G[�o�c�!y��]&�):d������OD��!�so�rK��+/�m������x��� WǱ̢"πf���0�PR�5Ā.��`u&z��k	r:��tG��5��B|����dC���4�z�m�w��������0~f�a��S<��F��Y�JT�:g�l�!���:zN�s�J۞/Y� X+��B�!�������C��v+t{Tc}E�PŒ�����A�Wl�S ��d�/��QnS��т�8��͐�G�iӑG�pu~�W��x����b��UPU�]����)�%	�p(ū�,�ՌH ��C+ѝ8p>��éa:{$' �aY|g��r]Ȓ
k�B��U�w..#�[Xw� �Ú�U�-�NGh�+3$�E��"��_�;?V� s��X��n{��8�p�k��*���:���G���F�%�R??!�ݟ���Pg��[����ĉ��~u�F7�ڒR��>�X�`�Ib�EP#��YU�6�V6l����8�39����n��J}^>|����U�� a�Z���Bi�GzeY���׮�ǳKp��3Kt�<�v�)�,�B�Ʌ�@F���P��K�f\����݃�d�j���VIH�S��E��,��VL���� +"Mr��V{����"�]��Q����h��D�� ̕�s-�=��_���9�����G"�aqO�=��D*h*p!���3����(V�����"����*����>���u�Gc��"� TQ�>8�1E-��z -� �z~���M38�c��,:�c�R�!�*w�_�E��t�=Q�+����#��g�6~;
�G���%FD�}=��O�vz�J��pa�G�,��N(1a"Å��fo�GY��8��Oi3��S�,�nm��S8��
L9�Z18ݻ��+�NbH��S��0�ϧ�F^V��ׁ�Fhp��,jJS-�h$]Tpv�LF��U���׻������FE�l�|/��4�o���{!ނ��|��SO�z��z����!����R��0���<����^ZE���ݱl�
Ci��7��#׸��?��3B��J ���de��j��I��q�|�R�S9W��I�:�F��h�p�eQ��`�dmXr�NOՌH�Ҏ��9�������&<�^辮�9��a�M4.2�ԓ\TC����Z��BO��P���D9�_8ye��MMBS��$i��)E���b�A��K�f��3U��l�5�i��3Gu��Xo�yy#uG'�ѥ�Mo^�%XcDu�C��'*k))[��v�Gt$�:���h���y�.�'L��Rҿ�o����Դu�P�:�E�χ��N����"Y(�-d��f_���sNg���)��s��uX�
~f�>
E¦��[��Ϧ��� �Ď-��U�)����.y!Ǿ!��s�"��f�Ⱥ}C�ͅZ+Յ2��2��9B��
4���J��YF��Q8ڟ7\��'9�פ@�m9ܚ���l���B���~�)��-^��
�= V�OVB�4�2����]�W\o�qPq��UX��e���h�(��]d���V��b�xI<A:q�@`$�[/�/�gV�G1���)n����ГU��gw6�S7r����7�,,$�YJPXtӪ;�0�8�43Yp���c�=g���nTc�9��{�@_�8���o��n��%�m��v+WWL��l�߮�0����H���݅8*��Jb1�a����,�3UsA�A	s�80���Iʁ�W��JLl8͊ > ?�ٺ+�q-Y��ё�Bx�yJ�Gv���F�P��[��*�C����Q�o9��K�h�Y �z����<VxY�b��@?c��~���L{C���a&��Ye��Wr]!O�o$=A��ڊW�1�숬\������^B�>�r�o�����EZ���z���տjfɗ�eG��r��n���t�����u��*����d����;v��8Ǽ�q~^I[�� H�^쁬I��6� _�ל����_Jl�gR-�l�w[!Ý�6d���6���E:&!X�XN堽�s��VWڀ�=w��nݤ ���f��4��D�	�v��������&���LUv8�-�0H �B��
W��ȴ�w�y�&��~���u�IK��6
�a�A�f�����3X��8S��a�o0�S�������/���J����u�>)?{���z!D(�w��o���#�xc�Z��˔ ��2��8��{�W=F
��*�.�:�Զϥ&�Vy{l��sMR����ϥ2���(�zn�����H����h�~A���Ezw�"���,��?J=��*�9��p��=��ɕ}�e�i]��n���:�)��+}>��>�[g������a<�'"��`U2��/
�yoB��B<��9�!������kr\�۷J �%މHT�?��������M,q{3՛[����U}���'l%K3��ٽ��0�%s`8�nǗ��:��I�\��Sfxpϩ��?�NbTж: V������E�j~c����+�c��D�Xѩ��.E�����k��G����	����L)s8��"��٨��C��:�kd%��}u�H�l�����aH���ε�����J��o�i5]Ij����F�I��a��Jq\{�-�@B�Cx��4�;f��=X��k�؁:��*�q�hHd�'��݉ŕ;7�¾��	 NA�$Z>ck�h<�-fjd��)�����������uP_���8�.-�l �9U5��"�VӘ��U�b6�$0��[��9�3!�7���G9}be6�YE��{�8r�����xw�*:J�Ț-��(3q�	� ���-��Ri�C .��M�^��;��Ci�`�xX}�P\n���9���}����L�$h"�>�a\t}�ʀ�p��e~X���s�T�u��~�D>�bז��Jt��E  S�6���+�C��oZJ��Ѳ�;
�ض0�X~���������Tp��Χ�Tk[�xh���3�׭����ӿ���+
> /�M����z��l�/�r� �=�j���9��d�.���YS�0��IQɜ���6>�?���\{�q��NG'��/��|��g�{c�[�Xyǵ�և������K�SV�R@iz�������:g3�-0p��2��a&j�14>~��3��o,>|�����T����_]
�r$NB����L �K$
��`:��Ԣ��ޚ�,ޑ����)��ա�m�Dz�����6�'�������K�c�?�k���J��
���l�묄��E[�^
eCz&q���6�S�v~F~�����OM$;�Ҝ�ֿ�`Iy�KM�� ��3?�K�J��ľ�f��N�Ս?01]JaG�.(A�J�����
�p���Ԁ5�CU�o���;�eG�x��E��־�]���}�[҉���x�
.W����q�&�I�r��&;S��=���Y��[�%�h��p�9���$��#Ss�)h����{� ][ԃ�+�-Fg��EN~O��}k��3��6���ׇ�5߃�k�l���M�sE�A�܃`�0p �����l���
*��M���B��J��F�}y-�QE�
�b��0��x *%Ƭ��q��lM#Pp.F���h��R�8V�8{�b��d�:�(��!� �v���˻��O���2"�$�3ez���ݑ��!^}�\|C�C�phHj�i�L��-�ڼ�ye���T��d8��%�螽��]uk�6(w?{'rJ�\��B!�~��M~tI� }j��.��@�8�B�m�����%��w�+07��.zj���;�� Xw�*�\�\��6QA����ZEO�d�
�h��0l��c��)��S  ���re�����i�pG�0J/.|�,d�W���l��i�#z/Cˀ�*�x�5w�1@ଲ�����&�Up�����Õb���S݃x���>��_*��7�-���:��b�,@��z`e���Dyj�50r"&ݭs�E���ܕ'-�ᑌ�w!D8|̜U����$���"��>��\"��mq����J�-��H��c��fǡd��������b6:g�*���ŋ�[�	E���,U��2����I���{�G�C����TL�u�m�f^�[�8������OG�&�D��᠄���E�1�	"��3�@9dR��Q�,/(��$gb����ȏ0���G�勍ǁ��Y��Zr�o��Ħ���I�kI�d$�ln��ٸv��k5�M�����v9�/
x)�����.��g�[p7�]ɖ�Ó7���ȗ�W��JI؈��xF��Đ?��%Z���{�I���E��|"�г�[q�x��⫐`�8q=�M��R�x]�
��V����O=#Y(C�Ry�w!�����cV��������p���M�黰9�"|AIڿ���i�,F��"��`
c����o�8�G8��=��������_�V^�?�Kw��ݱ�)�=6׉�A�������s
h�'��tx���`���%"��	��T�oF�{����y�L�^��9,��z�[����M^ �G��Ѿ�P�8�9��+��4���Sx��"σ3���,#��~�H4&���FH�X�M�סl{\A����Rn���S^Fv��`h������7��nr��b�G�|�/3;�����,MR%�EB0�w?�F� �7�ʷ�	3P8�a���A����ctj��H�礼��h�m~�����D����7�tƿ/|v۴"[Mc��ǎrL��> ���
A�� �%]z�C�=���a�%��-��%@+Ȯ!�Gښ����{��~IB0�7"�����j$y4"�#�ȿ<g&^�{�"��D���A��(��Df���c��Huܔ�x_�n�U��s/vC��Ғ�-Ux+<�B�Y9��GE~���x_7�%�+�`yBv�@Y<�2�FY�m�o3��F.1���5�+�/���*�tA�?ȶt��4*'�� 0�T##�^�W��1�b3_���sT�bE��Ğ)��O��2�X�pZ��0Yf�����g�;�X��:�Ԝ�ZvXq���q{���/���h�$�����Lw��>Sx\�H�Q�y�Q˗� �!/(�A%���~n��2�{ kb��J��y޳�6@]� Bz��Ng�L��O�63��&���╌ԧ�נq��)Ycє�*f"�6�)��n��	�V�E0�抲�o?��4|Zb��B7UQP�qqE'�͋6U�|�N�:�cvB�<>F�w�
KQ��
]e�\�#*{Iћ��T�:��hݣUe��:�4�t�|���f��HY8���V�h��Ѫ���y�ɺ���VC/��ڛR	��S$FI����oe�Xy�o�rEK���n*��1<�{����_���t����tY�P�wp�S�%�>+�۪��&��`~��t�j pe�������{��������ߴ�COȌCV��J��<��[����=Ku2���d�7�GpL&�>��X�ˮ�':��Ǥ�ǵ�2�"C����F2/;B,7�2�9�Ɲ�B0�3j�R�����x�ނ	f��Ǘ��N���\
��@���<p����%B���Z*�_ay"�qq���D�<%!VY�n<��fQ�\���67o�xM��o�;�(~y��^X��������,$�>��nX�Oňz�����A�}�k^�n�"c`!��д��������e9<Ԋ�N�k��G~%�@��by.�r!2~�]+�ᅗmm��~&�ϫ�T��0=~TVa@ڽ�֊��A���,i�e�Wrǭ?�;��7.2�ݯ���Y�43�����#G���[���`��>�(��YT�}v����B�[���~��tC��1۝�a�e�0&L���ܟi�޵P��-GUN��������f�^��4����;ȧ�T���?��G��3Y���b7u���E�5�������fЛ~�A;Wz˸�C� TW����� ��#�S
*�z/ݤ���I�w�Q4*���]�?T�����F=h���\�.� ��[�<�d�~�Ds�wh���	߿Z��/\����L���"/����>�e|��5OZQ�,f�K�G�<�T<f���r��N|�+�%.�ϰ�Iև�I��R�X)Ś���/.��P��a۝/
E:|���f���=��@j���kG�0�1����)4j�M�8�-�yi��0�U�1�G��V�n�x]w��r���sȡ��,��!�1�%&�$��h���5m��k��6��Yy��h�G�z n�%��R�c�IM��[��V��$�o��,c��(lu���{��y�g�K���.�E�-.d8�;;D�=+c��z!�\sei�S��릏i/���h�[APx��|�5����i=�%��f~�ݕ)1	��r[��Q˨�͔��#]-�NE�rE<yy����u8�ߴG�ᘌz0�k�s�8"4��ͷ��Zo��7W7�AL��L�ُ��-�M�i!Rے�K���~+q�sR�Յ�F�M(��g `��t^n�%ێ�1I��PF�����s��^��1��ĞL�|�ʊ��j]���#��:ր���l� ��K������K�Zj�쪷_[H���+;��䏁k��bI��T�t�%K�	~��!�����#����3
�:P�U����UҶ��䌥M�;����(͡]�E�΍UqOH�ڍ
ڥ}"�����w�x�����=���c��My'ω�"�gaBr}-�f�'��P���Wh7�B.����{��)����v����]�Wsnz$[�Tv�־K­��ЌV$��7g8��XΎ�R2{�o�X�t؝�YG����� ��O��(/�b��3�I>�
�s	EW��ҤS�9as/R���fUW������t�P�C�5���u{g��)ʂ�N�*����b��?�;�^�gU�QC�m�4j�o�1����5|3x=�x���>����R[;�R]l�g|w��Ҵ,ېr�	{*Z�5{L�����Hܛ��<��P�o��h&������H�+Ӕ�ƴDp������|G�6F��X!�t�I� �I}�}qT]��SS������>�ה��7Z�7ܩ��!��eOr��&٣>�ݲ�zE
��c_H�G�f(�Y�d����3����=s�� �#����tG#�ma�p>����B��l �8[(a�R�o����D��������R���b�ڍ6A�s��EST4�&$�$D\���?��q�ą�ϼM���r&?��[�^��x1�,�θ�U��r>Oo�f���`I�rT��ٵ9�%��6
�,�	�A&�m���0���ʥ�qZ�:���Ҁ#t���A�"��,H�	�m,AY�MP����gȐ������ݹ/�A�a�զ��o�J�OG��y���p��[D$�0�K���}3i�x5da�����ֹ�B��BE�\޸e��xm׳`�a�l��(����o�9�b���IG��웙���Ò\
@����P�ի2� �Pųu���ZAQQ����<�"W�!��0�֖R��<�N���遲�G�n@��ܮXiv����n�g�����Y��)��_
Zp����q�؛�a���;#}#�۽͡�uM�^�!$sX$C��&�~�_8������X�.��m���m�~���ʎ0,fG��k@o$µI`"����Ѳ[l���􍱰�%1G��&,D
q+���ߖ��9V�з
�!jt�K9�Vl��l���oI�hou�6���ŚU�sY`~k�pyxk���Д��%K�)��QUxX;*�:B����% ��p"�_����P�@�j.�s����{y�y��)��Ƚk����e	�YP^�/�/r����E�����E4!�������e��S��d���C��2�}��G��x���n�@�!o��:����Ti��(��G+Q�5� ;E�q�����������S��)P<I�u�N�C�tZ�>�)9���]%�����	��s�	N����v{J���x�]ALZij�{��Č�UL�[j "��O��
'���^�C������F�v��UJ�1β�G��1j|�Pf�<���/�����'CU��"՚���qZ�Y�jۘe��j�=5ηZ���2(�³♹��-V]磩����@����F��%3@A��`�Q3T�p�'66�vE������1�<iпI{	���ĢJJ1G�n&�cC�ff�,Yڳ�a���yr&��p!b��\�)��6�����OA�*��Q2�X]��S�y[��k��엇k�D��0;W�-��`_%��LR�������L���oU#2�����u^~*�%��	�}G��LBn����-V�'0U�hX;�E���.��I�?�-�Z���P��fp�����).�П��h{sc��q�kjy�[ȡ��gho7�!�&��U��yF�G_p3��nv��Z��8w�7��y;y���G��2�w����-g8�uǴ�@]w��TdP��;kYs�YP�;�Q_��q�N��ê�����%��|��K9m(4Q�	e��Gr���*�����N��5�M�<Vt=-	��ޠ�]'�u���*������'�]�/���g
?����-a܏��(!�Kղ��6��j�<��hڵ��A��k�G�1�������>�3CK�B�V3�	��u��$�mZ!��R��u@(umT�\W���?5��劂��֢ �K-��1��v�Uh���R�0ˇ��1��ԁ�Z��8��ӏa������& �+�'F��A����	T~�|��9�����.����	_�7�n����rj� (C��v��T��Rh�\_ڙ� Zn��lG{���$P����K�����nP<��4H�������(��b��.�k̇�Y����<�Y�u��N��
�T��cf�x9RF���MB�����'��M��=?�7r�������،4;���^�;}���o�Ӣ�Q�7��2̖� ��0+�\������-J�X�PU��l|��� �7�MM֛��T����>���&F�xn�!1p�$�-��b��e�1A������I�z6[�M�D�����չ�o|Q�l����W�� ]� e\*���t3?��΁~6����R��� \�s��mJe傀kH������j���2{���h�Z8�Ԉ(nz�4x��/�&�@*�Ɋ���b�a.D�/YşG.��i�"Yq���DQ� ���90�88��[�
=H�'k��⇋V o����!I�!�9�{iLo~@Pm�ѸߊW�h?
Xt����?��i�pIV�.����-�FI�ʘ���c����8�ר?mr2�۷��Ez�,�!`'`C�_�b��U�{���,��W0'E��D�����Y宪��=�o,�x+T�0��v�i�q[Z�6#"�=��ŕ_wllDim��;׮��_���^0#��.�0����ҹ��p;�氕��}_��s��@
x�	w�G���Z5f��»1>���1�lt����n�~����_��͖:�Z�+2ޙ��s�i~Zs
~�4p),��"�Q����
�Y��1f��2,+rP�T�Ɉ���3��4J��랰}
Q��r�DO�nw]��q�Gb5T8�����|��V�9V�kx���P�������[�ܸ��}G�P�t�J�/�Ǐ��������-�p;�Ӟ!M4K�5�W�����ei�˹�LA��
a�>�dh������gD)<���v��|�l:�Wr7���"æ�8D���c��ϴb�Ԉu�?^�}\�7��P{%���eއ�@��	"��عL�@�!����)
ٱ��r
��Yn
8|�zv��_���U��_��1�'w��D�1�vy%�qc���'!�� t�޴U���I�c�S�nx��ke�9;�R���AS㊗��}T�9�}��&�߫&�5�G0U�^�Y��@�k�$�H^#����5|C��Qg U�A~�#�(q#�H=u@�~��'* ���$=Ge���a�h�U?b#���z ���˹�O+��zQ���Ď)PA��J���{$aW \��ugl[�щ�.&,}Sp(�,%;�̇���h���%ܝ[h';����ϯv#ޠ�g�O:� &�rm��{a�@ϑmM����<��"�s��+ �/������.T�;=���*Ď��	�"�k�[X<��-Bm��||A�8����5�U&�uj~��3ϯ`a��D��縘�pѬ6J]���L��*ۓ��[�@���?���L٢���=X{>k,��0|�ޤ�G�@�~�Ik��VK(�c��`��XO�� ��(ʝ7�*4��!T���ī$�J��Ie�F�7�o�Vʆ�3Gk��ov}�n,'��!��z���ہA�
o�Pj�7Q�h�`B���:� -ы��2��15t0W����=��k��$�ckU;E��V���zrK���*��B1"����P|A�~Ҙ��g�٥��G�y_��M�œw�UD3�I�O$�g����d����]T�YV(�0���_l��f�R>'�wҨ��W�G��l������Q���]�є���u�Z5��ƌ!j? �ȁA����	F4щcd����G�2�[�fjA��m��j�jߥ�$������l�� ����\Q�&��o��,�����_]G�x]"wM�x�qw���y�Β-l���s�ǋD��BXF,V��{z41G�
��{��#��B�cB$��ع�媢
~���bʬw������ �<M�����JE#E�̢��)��۞��ߡ�҆�5�X]��Wb�a���.P�(Y:~�Tר�H�zɛ)7�E��y/f�F�D≓�q]!p�Ht����3�����>����߼*�6��\�B���fXc#r�	r:�х+ ���}&�����aR�Yo͵A�����2�;��;�.�[�B��wp��
��ݚ�6j�x�q�K:4���>��������/ڟ:��%�#i�I4Z��)�X5�1D��+F��(Q�n�z[�s���{�6��Q�k��f�5�X��4NJA����B�%��0�b���-��䯤wa�4�Lw葙�RI���W���# ����'[�1�"�YB�C���C���l̉8V)NXb�9��.��E�~r��
R[�U�9D�t6��R�����܀t[!�5	Ysn��%�ܣX��^�{Y=��fqJ�ȼ��!���4VRC"713
��#�ӽ"��Ǥ�I�����m�+A�0� Ў��{�n
��t^٥�.Ή�g M 8�(ju���ѩ]0*Bf�Y��E�����E,�e�,�/�4�^;H��t�D�2�%�(��^�\@����j��=���S��	�A�;����IpD�? /'^i��=`�N6�X�O>m)���IoB��A��֮6#��iZ&\����+�d��JKYtE�)_HT��
�0�0ł����X����/5�o�kYIEz��E!���a8LQ��;��"zk$h���ȣr�M�IX}�5,?�oNv�>J=�Cn�r�"���_�H�zu��5����0��?�P�J��Q[����oaa�:���iz���k�o���Tr�t�����B�$�av���W�ױ�kʜAA4�	�W��:W��e\*�Ћ4��ٰ{�����X_�ƒ��������*�ݴ�Fh���iP�����@���C�죤p�W�b��%��h7��'C��Q�	.�����v$/��F�È��FPY�������\LE�6$G|
�ٝ�Lm:0�� �{T�u�JfHi7�Nͺ\�t��IF�Y`b��ǩ��练�ZuQ���Y�88�i��@Ŵ���$A҄�>d���؏8l�_%3����`l�~*o��;勯���4#:+� ŷ��6@K��s�9�G�b+���6��������p.�$.L�iœlѮ T��{��?��xv����,���F��3�YA��G��?��\���g0�K��}�pl��ܚ�ݦ������E���6�>�^���1�6Dw�RՔ���
�0�t�qr�cս�io���[�a�c�L;~C������Ə#p!�k߱�5����[��j�d�G}<��!��|��*�<�#��aWy��%�W<T�������Y�ōk�G�\��xZ���V�b�3z�O�6,���w�VF��5b1>t�;qիkh:������"8���֟JECŏ��0k�5-��Aʡ:��m^f j��!+����g~�����+�3�`�'���_��|6�2';���ա�;	܈�nI����H6���v�"�@��3��,�=WiFr�W�r{�<�F!�5%����;H�A��%Δ����}*��2e�Ę�gy	�lWD�Lp���iK���r�	�L����&{���l�st��:c-�Bʅ���,���O�����~gXr�Fb�l&���}2N�0�|�p!* ��_�~��VK=�k��2ug�p�n�S]0�FT���<oW⇑+p���h���"9rʂ�3e�E��d�}�V 3�C�-�g������ڳ
o�5�r���t��DSbR�?YX9�`���F����(�����j3̐�5�%���` �o�1�1yx֗Ҵ;0�}���/����Z���*���\Logl��a�ϩ±7�{�.�d�C���q�(����K�p��/V�.0�E��]g�������	R"��{��=<\�3�qC��J��TZ��sm�)�a]�҅���@ �|?�x�5��R�*�ES�Z�����j�˭	m�|���@�C���v������,�غv�HT��ރ��)_�l�^ >X!�b�<��
1s�����{B��"ɀ��	�X5��)˕�!�"J���G�k��l��3'z�svd���X#��&G�N�ɻ"域��O~y��oևW%�=#�./PQX�:\/̬���@�=W��BD�?��u���W���Εsy���{ Q���7���p��ta�@�!��\4Q�к��ڻ��[��G����z�o1���>�VǬ�6�.xŦ�c2߱��uXFɘ��G�&�!{q	���Y���B��Sc�%a·OW�|X������e���L�le�pS����#:�SnM�>^͇��q H��3ݙ}�]�v�&�ӆ��Dd���r��*ZA'�~$�;l�7Ԇ,��3%3�k��y�np��/�[����=#՜n�-¹xv�� %J[�fA���<�q`�Ok���$^����9Е�q�U�����[��fG���墁�|(��"[�]K��<΂$	f��>o�Մ}��z�9�L, ��:��|8%
���G&xPyOG0�SUʈ�,�������@�sO3�ը��-�/IGi$o���#��B��eVP-���o]�v���ߙ���{%!Yt�ٹu@I����HO��2�STF���T��
Nse�Ҍ��R����\�K�/��{�"T+�p�����h�Q�r���0��- �J+93J�|�o�������#�ת'�⺼xD�O�t�
8k=���r3���:3��Zn;.t��QkL��]�h����v:���s:�}�'�����0=�.?쁽k��q���|�F ���1���*�� ��E�=�m 9a���&����2�����q$�Ju���8-�ƴ��m}��I�k=��(�D@���E��
R��;��Ά�S�A�NĢ)^׋,m"�Q[��u�B�6Y�f;�D϶���^6}@,����v�s���myl詅1;�TzK�!�X�1� 0���j�_��ss�xa����F�D,q��q���s/��kq��[nF�b7��S��~D.��p8��8�rf�D,���=�iŧ[�#��1>��<V��Mu+c�[��n6�uyo�VN�f�&OG�K�Oa�Ҭ4�P���)��쏋^ˇ�7�fI����SG��7{�g"���m��5��o��_.��K�#kx���(ǂ������+�N�>މ�>x�ժ����]��ޚS�ݮH�Ᏸ�����ڳ���t&��ʫY�n�s�KP9��i�]0'|�<�!M(�r��D��2p2�j�q�Z|�n�W�3MqвS��AP׋��vˁ��KSF�(���L8��6# �2��vippS�'_@w0iN�՜&Z���	��R}�f��Ҩo\
'b�N^i	d3��_1.jb�k��t��,X�
�y�0_)b+������X��~Wp� B�Iќ���G�my�x��m#z���G�"2���+M�
zV�1�N�V8��Da%sA9�gt����G*��l��1>��3#��[��V4y���8k��B�m8��x/��)hC�!��N�ͅ�j�ۚ��){�z����T�]��(�����=w�Au��s��z4�u��#���#Iu������K�j��/���.��I�7)m��M���ޅ����1�8�[�`F((�h�p�n���g�II6�@��)7�fg!�LoݦQ�w��_�3,wl2v�ܾG�j*��?��$4�*O}�������Ȁ��Rd�B�������K{(]���3_��9�Pv.sG��n7܌�?�1���T)�	�����.�7��8����rO]��u��j��w�{5z1�?�p_�ަ�b�](�s�1Rb����Z�P���l��9-��?�kF�+̣�Ј\���.\�5�b�M���Z�����t���~�f�/����LMP Q�E3?o{՞����*3���y���Fw{�pz�Z|��h��3p���z~^��*�̍�E��&�
sQ^�ah�h��5^F�#k�d�M��!����sw��^4�vP��ݑ}a��6|�:��`�?^��m�~l�I�,����p����;�69��d�8ZS�j���G�)��;$t^8�6�$뱢U�pm���l�E�-S�� f�Պ4� ��hr |֢iQ���a��V�������i��@��E=�_O�+2�R����>tdt��x�B�;K���}�	0��+��,9����H|��@We��l�i�`����O�w�!Y�i�f]�p� EP��!��2���=�,30��T3;������/��D��3O+�M��`�/9�6$�:�.����#TT^T?0�l3G���>G�\9=4,�z<���c�t2@]���-�1	�l��)�����{�B�Tr�3R$�O��5����`�|�R�Y�j�UC	��|B>@A�d?�ȓ��pSq��m�Y��.n	�I{~хi���[���������F�{$'`���]ut��H}���?*nOJ%��"IY�5��o�jPV�);"�,<|����k��[ �9�,[t��ugӐs�*�%<>=Nf�ӥ��~��/�?:�����1����	�Wi8������X`߾����zYS4���iK'X4T>�PHd8˕]c��˷�$�ڬ;���W�f����n� 1680ÛA�+ѻ(�u>��t�G)��j ��V2�S��o;RF]�eӛXr�C���wa7�W=�ɛ��Ё��+l�8��5�zsh>�5�ʯ��7s�����V�<����6E���Lᜆ��O/��:Vx��E��;���^� �8f4�1�K�f���꘠f�d@�wu��8�4�==��5�rk�.����A�&wR�㈟��� ��#�����K�C>D�m�{k�cDu����Xw�Z�F���*���aU)��ҿF�`n!�ч�d���|��ĩ�#D�p�߭ƥ��($���q���ɪ)n���t�-�iW����C`Z F����i={��e(�&�GQ�I��o�4n/�*��GV�Ǒr@�+���^l!�w��ԦT��Ay��{C����0J���Þ�\-�3z�zaڨOr�(l���P�Oc����?����G�S����`���ytB�t�4A���r��($��llA&	s��o��='XH��[�!f+0%9Pl��V�b�7r2$��97U���+�7t��\�ffl��-ɏ������+6e���_�2Оf	��ɬ��AZx�����g�8�[tÊ�5��;��1�®�C̎��*-NNܲe�����P���o�y�  �Q��s�E1�G���d'":(h��
׀�I��.T��]�����b���R��2�t��c<d�?H|�O�a~�z#�ѥ�a=[�:j��=b�"M 9�G|N���&&��cy�LK���
�ןE�JE��w�ڤ�5p����j�q��2Z�%n4"�����,�$�W�������S�
,��%$��V���^�jV������H2^�'���?��ߓ���{=�&�"2��CQ�N�A�h����̩$idAI&q\~CP$�D���|��姙�f���a1°0&ꙓ|&:��O!g��C��݋�"[}{QOQ��#%u���`YD�u9)���;]���]i+d�!O�q�l�tI_�>6cN�xw�M��9k�&��DW$U�T��>T��0�-��%�*B_��,��ܓ���J���A8~�[�N�m=Q��r4�T�܃#꠪d��WSL���]N��ipE�ɥae�	a���C=��є�S������ݴ���>��qu�ս�1n}�*���	��~��Ǐ��]�/V�ٱ��$<M��*��z�ֿP���������4S��Y��xq�S2ı��}&"��Xd�g�&��)+�h�0���ij�+4Q��v9o��1Nв�@��o�~jLu.�7��V���g�լ��m3Sԅ������'���G�X��j����ɨ�Z����L���ꏕ�l%DY���$�iD�y<[��w�T����Ӣ��9��~��쏹�����}�>@ZO ڻ�J��G��K�;�{���N�e17Lk��{�:ǩ���Wh�w�nZ�J!z��V2W1���B�s$�l��y��b�..X�jg 4������Ώ�N_�9���ph�D�}���H�^��C����ծ٩p�U���W�}�aH�R���z�G�ZO���pTwup�d�p�Jm7�3[W����DPh�Uϡ=~�Y	v�E���OFp��眏\G�D,�>[>�xd��9Q�0$�/i�ou�&�u��]��~Uld-���?r�� �|p�3J�2�pek�7��)Q����Ia�sk�㽡+:C���£af�����}��#��=�f��)O�Kd��7�i�������b\*��ρ����ӳ5������z;��r�k6~;�F7
4Ӫ��],����m�N���.�5�̠����m�O��-}U%�
��G���9g�'�-g(���x�m�d� {*~��L�r�I�ؽ�����n��:��ZyIE�W���@��.��)U�0�p�;TQ���>�ˊU���Y=>tܾ�P4W��D'ñ�0t=�d�:ɢ�\H��Q�Cȯ���sB9Ҳљ����x��[���ȟ�7+r���P�vNt[�D�^4C�M��[zU��L� ��%Fm쳃M;�����Ѳxp�?|8�T$�&3�Nfq��iUW�i�B�$�_C�8ȱ�`T {@\�=����_$Auf�.�r/�Z�v��?�>߹'�l�@_`u�g6�p�L?1Aգ���4]����K�2sr�p]���B��R��Ԭr�)%{���&��CD�f�srP~���y��"�fD2��������h��M'φ�q@	0^.n�\�V~f�����B���.aE�7�& �&����2 '�C�q�88b ��~g��p(j�{ؿ�[y�N>�mB��.�R�,#ҫ��G�CD:5��4>/�ԇ�������^�+�8��3J�D(�		�5�=��䇄xy��o{���s��
��$�k����Nֵ�Z��4f����xMrJ�J {92zT�d�2�j�S�,�M�H���˽�eJT�a�]�><��i�U�{r(�Wh����dR$�pv���� ����U��En}.�jmƧ�2����Hf~&��y��lĭ���Vd5�:�Ul?�d����0���٧&szx�`���KC��]��d�yW��Vap�0@r�#`B�2`�ߚ����'t͔C0Q� ��(W��FL�p��m��ۏ�+BV��$S���o�1��.�Ȧ-w���sFhPT3p�zx�&"�E\�u�KL�p���G*\��f@�N7�$;6]�E���/��] f�8�2��b�4u�B�:Y~V.s4,v����-�b�8���T�;�4�i)"��1D�+��+����g��]����)�W(�����L�0-iM�_��{����ac0�i�(�i��3��0l:EjzȰ�$���0նl�v���mI� lq�}"t�V/����j��쬧�δ`���A��s�bׇ��Nhb���ڬWcB	t �&Oc��G��+l)xR��0���V���.J>�sak	�*$�M*hhc&����"F=R}���YT���\�Ε�a�\��j�?�ͣ򃀒C��v��'�\U^��(�����6�j+]W�^�z�af?}&���o���A�bQz�S
^u٣�w}���@@�Z�:�ѭ�!���X�g��<����3B�������jT&�OG�k��Ѓ=[����W�u)=��n�%��*!����J�"q��V��O�иػV�-�sg<���Vf����ׁ	R��L����^���sH�����b�Vd��4��4�wC"�2���+��,9��H�1�HQ=���/�~�,G������*���}rj���
^v����*9� ���'7���T�?������}-�����k=y�*���v;|ʺ@���mDLz;�}�������D�O�.�Q�ve�J|�֓@��c
����[�&��-S�c����hEr�<y�B_^5CɊqŭC��h����<��*t��n�$���bJ8�����=�֏�Y�i ��b�p9�����XY|l�ϕ� ��ʴ!*��K뙗Lp���.���ӝ:�kZ��*�c-��q(V8 dhK���5�񺦋�ш���ܔ�B����A��4�6^g��7�5��l�.���[�:��&��õ��|�+�Ef;q�jj��9-Q�)�a�����:�*�1wck�ӊ�"b�UU�܂��=���o�l�"M�1S�2~��$��U�\O���wa��!Qn�a{/Tu������z�F� |�f5Uz�6�:v��<�-�j#�(!�X�L�e���ܲ$ͧ{�����=������M.i��η��TG`�7��##�F%�A{�q���o�Q��P׮c��d��"aH2*G/�B��U�gZ�|������JA��)#dcp%�pY��ߟ��E7@�͸���<f�rY�5^����Z��J^�*�7ܸ����Et���:W?UN����>ȘJ�e|�^3��
?�����(�BY�������(D��@�Ѷ�9�%���M���	�}�Z��
/����#V�ZCa 9�qQQW����4�Q�/��OМV�ϗ*�;�ϻ@mYQ3��U��H*� Uv���E�n����" 0�����} Aj���Z}�ɺ�=��/jآ7��)��t'i��ϳ���,�Č�i�Z�p%D��n�/T�� �q���i6ه�����	q
�ܠ^3Z��2Y��H���t��Ţ��w�6�,5�
:d@ ��I2:���{��h�Ż���H��_��ߣ� M��GL��\>���ST�����y���t�r�]2C`�5
�A��2Fu'Y���`��̷��$朘Ӫ3�xc��$^�^�7�qYÿ����
~p=`����C�Pz�s(��s	"F��F�br�����P���e8>�.d���v�d�HrQ�QO�>d^d|��c�G���^"��st�,���&o�溄5�t� ��}�O�����b�(�QP"���� 6��j�9Ch�������?�o���+~-�Y�l���4�Y�����'y�J(�ߺ,u�����-�f��(����x]��JV�&�[��2H���vu��f�����v�5�,��U7� �����̤]��'��3�Z*lˬ�||GK>��g�.� (�����,�H\2�� dWm���e����w�%O	�"h<l�ئ�k���J�:��^����)u�"$��3oV��"��3��8��>s��gel�,�q�#��3���s>�Bmb0�9��������k/�645u:'rwԆ���"�BN��z������5�=Xx����yt��>�C�<*��,D&S~���sf[*�1,oաܛ=���y&r���;���L}dYQ[{���V����j������u�߃-h�u(������9J]��5֡�:����q���JX]�n��K�1f8(GI����O/�q��'W��&SOV��E�l�"	�o�k��mz�$��!����eU��U�P�>~�7���y�֋!&>4iq�Xҽ���uJ��#l&�	=��߯� ���^��|oU�"��߻�����5y���-9�[J8-�.e�W/��-���y�2�T�,��),�
L� �s0tXǟQ���[Qh��Y@y�3p!]&@��A�3{l
v�!�1���cb��S9cv�L�?^1VD���M�>sڵ��i��'-j��1	>5u����:u^O�"fd�e-@��� n���Æ}����g�OϽąy,��S�s�b�{M�ϵZ���7��[�N�!��$��s_C�~гMa�^Y 9F�q����&��졑~��j��?���i#�k���b�t$aWI���ިa�G�#�T�>UG-6��������{�m3M��J�� �D��P���Ǌ�5���9|���*�\"�90�\N��%�=�ぐC���˅A���׋R��f��6$��fo^���c&��AQ8ҐA�����_�Cm2����5/O~�/!S���\VCV�s�[�V8�b!��4aK[�E(�_�|�p���	%����"�W{.Vz/�<A��N��. �Kq�h���!��U��!c?1r�*���q�x|*��i�"����ڠ��[��&Xl2�� ��|�U131��u��W}�yx�D�g�Q�Fq7���[+�����i��o�ϟr��kW �O�շڰ����-Esz<
�2��){��'��-u�}�0�Z�#�0ߟ|�O��V>�P�4*�ñ�`�gP�k��A�!���D2D�P����Ė4C5>�qd�x�䄪m��\	kC6��B���%����Ɍ}
~x�#}��[, ��x|UB>�A��i�'��D-��&�f+X`�d�kȡ��p�@�3s�5v]qm�����/�X�����kuqX�&X�[��L��Q\a@`���m�Ud-?�K��".^x-cu?c�n�e�����d:=�ғg/=܃be�	*+��B����)�bT���(?�Dב1|�|����sPCՠ��I��sX�)��Ŏ�O��U��^���x(���E<8c��y&%�i�� �����eHs	�ʨ=������>S�l"L�*Bf�騔L�Q����^���j���1G�Gp��q7�I��9����~G�zv	�61��b�,6T��Bvw��������2.F`@�!�KA�������84o��9���Ȋ�,�yڭ��I�<@Q{nDF�zx���N
!�K��I��)ô��LQ�0d[?���C[�t̍��r����Bh�"�{����q+�V�Cʦ��s76��ƕ�<� ���L"�#��7u4OA͝��`N,a�{�鶌�ji�-G��g�Fr��`�.9�s�]Մϼ����)@]�0�Js��9s�0����mr��������?=��ϱ#�#�䧻�s9��}/�(H�t���L̴����gR��4W	��$u�&n��c<�"z`��JZ|>vܢ�/,vzZZ�-��_�Nɭ@�!��^��L���L��G:��H ,�e~�̤
�h �A�O݉-h��j��s9d*��}�V�^qCY�pOJa���HyK�(�!�yQ�u<�Yu�X�Y$GĲQf]��n����p�/���&@M�������'*�Nd�p`{h{
�8���4�yP%�c�K����m�'�ʡ�L�#�Q��Ҝ�B`���b"�����^��v�X6I���|Mݸy���X�u�Y_�o��([�!�(�j�hd�2{�����蚝R�!����V:��ő"y�W'�pB�W�$�l�lt߀����k��I�#Ags��^�O����d��>=��n��:U�ٳ�_X�ep�1#���{��Wõ�?����c����H�n��[S�Z&H��٨/��^�X���G4���ב�S�h���[SSԙ���4�#a�\��x�9z��@A�z�GGz��Y���>r���Y��WF��p:n ܽ@1vf?�47��(��|��|�z��� x6�MsZsq�B�{�����n;%��C��x*�&gѩTJ��k`�4j �����F��|��촌�,ThU�|��'���O�i��:N4�4�̹O�mZ{�#���y 4�I�jZ���qQ�tY�ϓ׽�o���>�
Vq� �;�X��Bn>�{'�1"d�]����i���b��Z������엗T����3>]��h
��ʝ�� ��1�~� �V�g�8�a�9S�Y!W���j��5gaT�J���G}���G�A����U�F�cl�勬�����gk��yM�ߕ���;i ���u-8S�6�t�j5r�g��f��\)8�_�"�B[�%^B�QVa�DJ�f�쫁z��#`U�7Dkb��9��O�̜2د�����.Jn�B�@{]����պ�\�uRa)z|��f��aG#�~c�z��9��6si
?s��˘�á����	���@}����:����
OQ
q��%|@�֘E4ǣ��$���<U��==��>�=� �������V���@��-�Y�;C�v��`��O �(�r���_�|���a6�Q<H�S���q�|ý#ބK!z�
��Ek��NM1b�ʥ�ĞH��P2U@O�}j����6)����1qp�_~�;�6��Qs9yfI`�`�-<�;]��j�N���G1ñ�`����&IwJ���oV��6�a�W�?�YbIς� ��^EnE�\�|��A&P�.<0�ig�F&�6����t�~�8wO�s��I%�܍�φ'I�L��ޜ
m�����1QY����Y�������$Ε)����3��x�O8@�X{��Cp����M��?�� 4ϙ=H�]�r�Ŋņ���g�9/;)�#4�v�n�J�qm!]�o��ݟ�����q^�#T�y��d����Z����e�޻�}3���^�Z��x�l#�v�[<#]���T ����%�	�S��  ���p�1v�<4뵕� Ҧ�B?�����RM֯�L��n5ۦD�?��(���-�J��������I\J'�+V���ȑ9��Ol��;�	��T2�����6\Q�~��Վ;C�x3CG3��:���a�֦nC�/<ٜ�����P{z݆;G(�kIkm�T��\�	^��4
ѧ���<f��I�a�4R�/�����I��g���kΏFb��ה�N�QX�����M򧈭a)}��aC��bYB��	;:���g�g�P1��������-�<��d��=�_����(�9%!�����D���My{E9*���=g���]����.2�VT����3"����P�+��^i�U	"p?��Kx����AK���eW�Jos4���2"}����oՍj�c\f*���F� ��Q�f���g�! �8�6B�K�# b��sHѢ��[f�����<�}����!�n'�����)>3`]��y� )�(�7�g���w�����"l�m��8�8۝0���ۃ+�
�oK���8]c��%��~D�߰ǥ�:p�%W���pY�{��y4�!Y�f�W#�gk��1�QWPڋ�O+?}5�tPb�P�p���%��W���?r�\3j�S||��ifг6x�D���4�Hj&!��F�i��z(�O�f��c�l)�{4Q�&T!�N~��
���6�rs��%$P�S26���Op�١\�a�h�a���=����B+f���$�V� ȜJ`P o�Y����0K:a����r��H|JRp�!益s_���&�����&Z��h�P->��'�1������ܴ������3���f�H��D��P]r�"�7]��2!|v�S�^	vL7�����8���ի�����C�q����Te�P�_H�϶�ɠ�K�J�׸��	���;�v]I�� }��ҭ>vщkc�A��­̆НL'4�Cx1U��C�ҁ�1�@W�ؑ&��� �s�o1%=PL��ʸ�A�p�H�F?M��q�$��+�Y��A�J"6h�/Q��2� !�b�ԍݎ2��()BO�>lN釻Ƴ��-D������	!�V<+�R0ǥ���0��iV=�pnHp����%��slIjJ].۴Z����v�k���Rv(����4-�$��ט�����5�-���mD����-�5�m������)b�meR�������^��V�_�(hqE�̣߫Z7ᛒ7]����T2��H`Ԙ�����A����_��t��W&�ĭ�;�߹]�F˱��PS��2.����b��� 0�蛹��1.����KJ�v�J�d� �������9E�e��إy#=� �2v�Q��'�`Nҵ'_�GT�ThLH<	d�W�[�M�$Gz�9�`��^�N&���l���x���^l�YQ���$]�|޸/�����a�X�q�6����U�T����&Xxk���B�U(�<W����x����Lb�X���$)M`m��y ��u��N+H��b1A�.��Z���`kձM�_�_$ِ�!���8.L??��*�6�1��7�;�Y�#m�3R�]�����"�9t/�Q^��cE���%Gn���Ԙ�%��4.��4L��k��|�Ι:�/����J�7�jvuH~�sm�Po����r�P�߈ ^y8AI�Lt�)�Ib�!�َ�i�������(m���e������s����-V�d�ǵ�
�``˷咠@Te���׶0�w&�ԣ<S�H.����R{�C�&��w�*Y�ԩ}<sGj�dͳ�eV�}�p�2�����`LJΦ����V��ɜ���g�%�!��أpsLn��Vq�a�Ԑ:C�	�8��vf��٨[���J����h~��=q�ꎲ;K%<���Z!���M�dʌ��3l��f�~��YM�^x&�.�y�!X�B^��J�+Y�,ff�<��f�=���Xu /#����ig��9�L|��(ח�v3��x�VT=�E4\���q�~c���M�CؔJ�E�-R w�'�Fz����=gC�*۾�Y
����6���1!c*�H�'H�=��f꒷��A&�g�<�P?-�v�[J��cb@���N��e������}�掃@�C�wH�_  yT�\�"�Q��i�`1.�G<����\UĘ�#��]%��XtP���uG��8Ӵn g�\o�ǔ
����oy�N@bï	L�y}Z��gX��Wa '!Ի�H�<��8��y/����}O,�-�8F:�bBF�V�������zf[7�[����N�T I e�)t�v�_4lL�\FT�EK0P��� �W���dTV�s��W�a%��
��qX�A^G�WC�	U�F�?|'�<z�+��؛f��F�W��N6��
d��l�ѽT,�	d �E@����ԙ�C!P֦���>/����KY<�ewZ��#���-�l�% P"Me��dՙ.�b�5����I�D�ޫ�ZBY���ưSI=j�&H1��[D���jD��$.0�G��b
s����p���{7��YT֋q���@PN�;M���9���t��T~Й��� �a*�q�f���R���'S�[>8��ȇ���~l�5{ɯ�D���S+�e=j����,�n/������d���A��
���#;�+i�V�9P�ulp?���J������)��X:��9���}fZ;J]���c��NPʶ�&��''����)⹚��R�� ��	�8��Qs&R�'��TXc��{�iYͫ���6�?�$�����n�0t�����ܻ��7��@���Gu�hb
�mF�8����:TXn*�!��V�_����Ïpz ��5հ��[h!���9h�TWX���8�6���]A>H]�s�z��6�Т!���!J�I5�k,���bN��k�qs��uA�T���r��L���ދ����?�2)H�Aηy^n|��գFUY�&F9؀���� �,獿C���pq�\b�} �+A&	������(4eE�w�����6���i����^�%/��q\_&z��UY>A���P�g�� ���-D�R`��An�ivU�Y鳨x�"ukd��/�� ��LV�M�/��!���rz�,�wr���x蠪�؍�Ď�W ,S�ۯ�����A����[30+��^7��;C]#�Q�p����ɏ�%U�\����p��x���Fa�i�*�#տ.-��D�a6#�B[ �)S62S��/�M��a���X�7�+�� �>�BN碖�k�Jh]��UW�EXv��8�S�F؉1[_�>0G����b��~9���~g��L_-1�s����{P	~x�钒3��e)�d/�a��h#�(Y����m�ؐ/�����Ay����c@x}y��z����ZU��us\����I��~b/�p�*Vk�d��G=u���HГ��r*��0�n��b7���M2�&E��!TS0�)��%��H������,t,���/w3�dh�B�F /V�	V���x��a�饁g���-7˕9`'�p�/?��p�0{P�zb->���ɽ&���m_��>��w/���Cc�IL���<uT��
-��$A&\'�����0\r?�z��ʹ+��b�Ea������=S�K�$e�Fј�k
!��ް��:S5�zι+�qgLP�:l�U���V���h��a0�Ġ�'+l�tE  �����"i���4�f� ?ǿj���$VY���Gh|���U�q�aG;"t4 ����>�y�~�>����o�(�l3H{�80����X{����D}�6�Q��<���P<TÃl��)��-_��S�3B��ϼ�4_Q������T���$�<tV�J�,l���5��P���	v0j����Ҡs���]8�t#��Y�7��Z�"�pYG]"�n/�m4���>y�6MWc�;U����:rF�"��R�a�^]�����O|���
H��W���&�۵�%�g���D��ը�nE+km-&�q���?T;ɜ@��,�5H���]+a�x �É�cD)�v��"Y7��D��E�=1�b��I�Q��6�~t?T����HV/��W5�6�M*���$w��5��ȥ��#m=�V��tL�b�)�H��~:{ъa�VՃ�j5��lQ���a0�A��B*��0���Y%V8`l�hg��!�H^�
�\�z�(s1�t4�Y�:��=�g�����e�����/W�	��blf/L�=��ˢI<*�9v;|z4�R���ؼ�W�HS��ͳ������ȒHZe��*I��{�u16S�?�,�?��c|p�p��m�+B��S�ʬuC	�]�^PJhT���^�4��=(�]���dOk�!;zm�n�(AX>3!��P�l��-���J'1k�ͣh��_k���;D��U�o:<,xs��d�v����g�B˔5D8{\l[M'�/��nf����'g��H��ʞ���qn-9W6?��I�d����9�dw���oR�6щ�%p��5-ڐ�)�6�"tq�$�/�J��I��()�ovKѝ8����`B�!ܟ�Ik�ц9����>V6���ne��V�+�)����:�<�C�T�(5Wu�ͩLh��E"��=R�[�]��C�M�3�A��@[�W�x��˵bR� y���/Y��w╽`�HK1"���*�u��-�ORŖ�Bb�X���y�f�̞L7��D��t�^YrvN?��eT\f��j���,��PQ�~���y�n!�*�<"u���e}>��|��xR�!(�!FE�K�������;_�nna�g�.��A����6Y)���vg9��Wsl|���c�����>4$spOωqb��&�&��Ew��(
���(}E�h�=��/U�o�ݓ�r R�����f�z�m��oK>*U16$��ٳ˹�I��c����څ�;]�� f��%��R��r��_���@|�8ӈ�o�];�)�7�N��-����b(��eP'�ʆ�J�(��z����~�g��w�h�[-�U<�#jM�՞�<�3��-����T��ȼ���>�v�[W�1H��"�o�� �L�i�#7����'��%���7cq� ��r�q�F���e��X�&q ٰ�����������"�pg*����F�#+p�p��VO�ۋ���r�KE
����(J�P]�ر��{rj6Z���$,4Xc���l��1K����*Io�է�������J$:4nb��C��恸@���iN�_d� G�\X�|����6M�o9���u6��������Efe����NZ;Bݣ�����?i���~�����!�$���R���[x,�Ru����Jh J*��6:��M�G�4T���	�f�x~,ܩY��}N'�C���,߯e���F���6%�0Z����k^u��M�(�z���T������?�����-G*w.���u��@:�5pV9�dwn|u�Q�¢�b0��$�v�c��P?��}�������M="��,^�=�k����?�1�f�g!
g""��L��|�f?��i��H5|5%�OBXa�;�:��*b5�~l�_9�s~k[]�����}~�����1Z29x��-�(��G�v:�5��4���wcS��G^R0��9澗$m��E��@�T�U��C�P@-�:ډ]S� 9��a�����Z�����Iol4jc��<"p�@����,1����[=�d��:Ʒ(�[�|�)�E��$	��4���Z?h̖��_�O%���/�������{"�'d�ϯ�*Hw���B�Q����~a|�;� ��C�.g�H@j�Hy��r\��[��5��?�5����C��y~#� ~Q��e��?�m�����d�~�l���&n]���c��K*0���V=�Ig���*��Tf�:��3'����9�X��������a�^�����S��/�	����&F~Rt�4A�*8����fV°�^Y��o�F����W�$�\!�-e��x�@7�L�K9�Px1] ,��w��8��u� ܂ s��M.��,�R~Q�.�*�����;i����]�a��SX���!�ą�H����pp�cTrѭ8���y�>O��^ԏh.�}�yr�X�� ��5?���v���d���>Ժ.�/�������X1LʜYS#�R�)]Eǽ����P�mP�h�peժ�Ψp�\��ƍ����>;v3��t����������P�Z6�z���[�����p�������b���e��o��y` �&XҥX��*x�ay��㔉��O�gb�L��{3�{@��	�,wsw���TmTi���<@�͛�U�
���UWTD2��_�D�h��]�^��H@�����3���Sn�(@Hk3?da�>�j3�l���/M��=���v�W��=t�s�pJ���|y��炇��K>���4x+c�2���a^,g�u�cs�~�Y ������4g(��gF���RA�h�2�_0H�-d�-%y�9���6K��1�C�"�d���*� Xt�:U-s�OLy�f��2��t#\H_��%4d-=��/G���e>���e0AL��,X��*�5螵�of������&F��؉�&��WD�h+����s{�J���T4�~��qIc@0K��r!.�}�q�V�̎���ʰKp�� Y�7hŘ�Yt�U�w��g�s.��>��̦-ڏ_:�V�JU�mW=99^p&�<P����[Ͽ]�R���C�����.��4��
 �6d<�Pk��sa}��f�+�nYn��Q�r�~�M*��l,�k�
�$�P�dש���'e�y��1��<���]��"�NP�[��,^�GQD���{Ǘ����\U���lPԛl�Wiθz�$A>g����!��S�Z2��;o�6;;ǣ:��7N<5`m�v���;�6�}0��r#��<��ǋf��^�ڜzb��}Qǻ�o|�>���{L��=����t���'��0��v�T4?�����q� 1uJH�v�*/i��k�8����G��Wܸ��i�d�9��X`��njd��Ѹ�S�~ ߵ�{F �3ESr��Z�W��%��m�j��eh �@$����]��
�q����	"�R.-H���} �x�qb_%��t�ٟ�-]�g��>b��F]����S�=��� ̌�O����+t�H�+�W��QQ���� `8��s�u�X�U�=hLC�u|���P��ҖN��)^��C������4d��g�B
ų�Y��BY��_�e��~	y_�1BHp�$6 	5��p�u��P�g�kZje��D��ù*��]()�+�;Y!%uc�X����|V<K.C�JY�{�(h�سJ�`�i�ʯ�UH� ���:K�"�Cd��.�/��O��ծ5���~�ѷ� ݓ���������'p(h��O���*��	3�5;��ZSD������3Ž���8P�7���r@�)4������S�1��@u�<�[�t��b�v��e��
1((�U�Q��?���" �'��d����D����xs�}t(����L���]����!p�)��F ��UÏ;�����-*�72B�2���_ �KM����S�?��L�K�����l�qØb�h�MZ�U�#��"^�+�@�/~�+�F[����RHK��.x� �����D���نmȠ�AU��"l�����.��9�ZAt���`��L�	2�?k��k��"�bnC%��� 㡦�
����s5s<�4�M���1��/@i���],�M�,�u�c��ܝf�����u4�Մ�U[~������<�l7zJ��a'
���s���Z`墛>5E��~F��7�°��6��i�7n�Gs��R>R���&D�p�_�}�!���p�k��!��	�O�-꺞�#���z������4�"��x�%ilP�y"%׌wQ��/��!{	ed1�`"K����q%Q`�ݠ��y���ǲ��jm���|��m��,v�s��w@���G����d��S[���s:�!%7�
�sD��o�k����g�f
HR��X���M�/XB��R76�ٿ�l8C0�[4�(��z3ayoM�;}�x�,%�j:-�g�,UN�;����{R�r��K^�g�#��?�/�C�8h{|ʾ0��t�L9�A��W�zI6��
"�}�*T�����͌y홐����K����Xb;�Ilhh�)��"1��[#!V���;�b���l%������R0����yB��<ґ1���pz�Z�խE���\���eU$��]���ܴzc��X�YDw�9/ʇ�;6Eg>��OoAJ]�J��<������'��6R�G9>��:oK:��.��q�b�N����(\G�T�l!��>�5�H�� Z�L���ٞ�w�����N���&�Q@ ?׽�"%*�=X�
�p��	c���+^��߈]1$0���F��)��,B���@�Fb�G1�����Y�I���c��Pw�`R���s� :�8 �"��	�ġh���t@�ڇ��J�wv&8%s�u���Y� ���N�Vr��=C��s��9��2?���q.��Ǹ���6 �k\�<7[��=���o�%z��F�V��}��*.?b[��2�wBVX�Z�} ~�,OU��\���TN�/�T: z�^��$nY����SXf�e�}*ĬH��yoN�r.o�.�~�8|���S�'����
�m��0Eq��ry=�e�̥5!Юg�r���m�/ԥ?	[�¸<����n0Y),�>�zK{�}��C�2"���(r�zj�5�\9w��� hv���OS�0gN[1�q.a��y��ԥ�Ȯ�W-��-����RUơ���+F�K����Ve�o�"Ԝ�J�XG
/z �/��J��ܯ�E\��a�;�w���NIR�EA!���l�RN�`spT�k��3�^�k	�\�>��伕Q!56�7����DV6�M%�/���uo+��#^�P{�ߋ�D.ð�z�\  ��̑��-��R�AP�S@�/�>�%�Uڜ᜼k�yM>�/�B�{������I����$B�q�9a9�y�"����8��#'����t�<w�偻y��|?��7#���x��پ�w�2� R4cX�v~꭮������C�ߥ/6��L`�M3>��o��YJ7xu	i�*𤡹Θ��"61�G��񯷞(����mu�+f9�JM+��u��asp4��O��\�7�pi�K�w~��_q�b_|CY*�ײ'�G?{�*�%֘I4�;]�����9�V镺��:jlP��t�������\���N
��]x�4H�y�.1U>�����{�I�oD��5�؆��>�g��\�n�j	lꁶ 	�w�@���`��U�Qo���'}��'�y =���SBLr7o}l�YbV�����U'�
ԈN��(?fqG )����=՛���ÖS�gy�_}�gx奥Q�FֶB�^�\��Ԑ�_��V�����-�1{�Y��'�v�U��늸�t�g�*���8��^C%�#��ex� ��R�ɕ!à���]*o�M����,���=/��eI��헼ަ�����.���p�i��:�dp�h�Ŭ�o��+0񄯐��n�lJ��E�:�5����2�w�m��� ��Z7�1hX�����o�.��`[;r�W�﫾�+��=�&!�iw���� ��o־g�xp�z���\�FE^���R���Z���^�Z�q
�2Է�wv<�H�����+��0���P`����e����;�h�����0xh��U�h��E°��9�⭵e����!��FR�l�A-�a��1��G�l��_sH9$�1��&�+^!,��t�Rϋ�1�\A�81���쮘�{z$a1�����(��þE����;�� �"��zҡ*o����.囃�]<	]�`�2?���� ��o#�%z�l�JmՍ#��۸�/N��͗/��bS�)踏/�����c�]���b����������e�R#�C���H8���x�$���37�g���o��|{�*F�09pi�G#�(P�#�33�H�8)f�G�S&J:��^o�5�v�W��-^ �EL-�IR��"����Q=�Ϝ���@���H0�-䮄+xwD��L~Z�Go�AU�]���6=5ߖc�^lJ(��e�8�HFOE��8��Kg�vO	р8ȏP_�-H"�Qڥ����t ���D:^I����3��g2,�P��ю���(�g�ShN��U�Tm�?0
d��m�F�OުWI�/�ǈn��	�ZM�Ks_��gGV�a�;��ܖ�!�:�zg�td��S�y�Hz$ꮙ@6�&����г������ę�^��4yOD��2j�O�o�,.|����J���V��a��aY3��4�h�XS|�o(VfGK��[?���k������Y���.3��Լ�}��w��v�z�t�o�84�;0ĳ\H�W��%���
�/��6�>����cw��*�{����l(?�׭�h���h�+̓��l���D�r�V�Iئ��q4� �����
�I�5F&x�0�4N�Z���Xc��h0��-��u�qb�8I�bO���#�K-<[9R��m{#c꾟r��Κ�۝u�9�����T�%p�2pWR�hԣX�B���f��4��Cs4l�y��{证�Ht���:��KJs������Yb�Zz�Kkk~�k	7;�7�r��|8%�f9,�Z8n��(�,ݒ�C#��[�s�����
��鍱�{&�N$F=X]�ܸ*3��7F�`̪���vT'Y ��;a�@̣o1@�����3� N1�
VL�d]�/x�@_�kW�;�7=2�E�35�-�3oZ��T�| H���'�OY�lp�۳0!��:6�JO����l$���׵�u����B�	#O���O#8�M�L)I��C;U��70��2 ��ɏ�)@S�4���L����$�b��O T�˘�����x�~"9�u���
XK�{��"\��)�u90�C�v=��7��E�|�&��bvӛ�� �a
du;��"��*6X�d�<�ML#�?8��_]掛tiu�%��(A��Q�Z��|sy��݂5id�Zp�FD�gK�*�.���У������$�A�}�U �����X���22���=�����ǥW��<>��b��invm��[�>[�&���P��~T�v�L��*���"A���Xy�d��
}��,�a�I���Ye�Ǡ�J���;��nz�RJ�D1hs����:>T�C��.6�1��D��r
�!ܜ&�'u�1P�p�R{@���Q�y$�d���{�_� 찀=A�"F��o�*ք���r�/Ң4��Ű��S[]��	%v��ɓ�5r��r�n��^�k�g�q���5���Y�-_����)Ufޖ�vqS�7tJ�D
���D�ѫ��B́��cc{�`�$hI7B�}�����毫�D�p��'LE@JY6�u.q�)����7|1�f!�H�
\�c��אl*x8�_X���Zp��P�s}���.�gG6O��s��l���\9ɜ�hZ,7�2v�#���oL������JتG����_�\��Y4���m��3�J�j�łP����V�5M��oLl8�C$�2H����澛�rz�8K\�r_���F�`r(?�+hȷ1����z]L�3��.A��]����U��˨����6���d
� �����!��d�ɱ���3���� R�Y�ۙ��g��f���8Q�Z��*\JL���
��7�s�%�0Q\��}���XI�*ܘ|LLv0��Rs��=�c������IRӃmrd�1E-��]���V�L�pjA��"o��.E�x\$#4�T|�e	|w�@������X�c�B�tXp	y�ՊS�2]M�Q��[��ȑ��9�<eTҪC��a5<=�䗛���W �w���)~0]��
�(�v���������r�׬�I������[��SkM���� ^<�1�R$&�:v�;f��<�|l�Ђ3>$��'�6]v�����E��Ɣ�\ }����g�iLFvَ�םRa�(��y��9Y�e�-�S�s����К�-�sO7�5�!�b:��`�'0ǫ����CIK��gh�qQl��CP�/-͒�Rt����I�9�C�*G[�.����5p�b�Ֆ���1�̮}-�oN�~����$�Y������ٓ����q������e4H�(��T��7�=��M�L���0Ɠj%uT.F��+�a)J�@�t"4��"�& V��+?HE�Z����`��$����n����$��9إ>$aV2�A>>[�xe�I�����Bs��o���M��q�H��b���E������c������+oy��*��|0&�筑b�"W�a�ҨFj8�{��`�4��Q�^�Cd@��l�
�q�z+;jZoy��PY���X�A�oQM4Ѝx���)�}s�K櫦��ʏh�Jx���K���zO����U�7���t�\�NşV����Y�䪋Q�}wfg���A����3˰�Yk�AL��\s	� �m���3�����t�=�x�	��+_v�>��51����X`�vYi��u΅���(Z�A���u|@�V�v���O-�<L�]��`��}����93��6�W���ڬ��a���襎�w��wqA������O>1��z�t� �������r ��\�B2◲15:�0����_��if��B!9h��A�L�#�ؔ����"�9�A�6� n�6<R�%B��F�l���H�ɭ&�?��K�Ъ%��4SU�L�CV�?�aO��'Cߊu�EiMΏB)7Ua}�U�<fn*��������Y��ʮ0�J��y�x�����1���ڹ�#�A�^_fiuM3T���"�Ml��Jo�C1�El�Z�f���=���s���(�@���h��֒��1�ǢR	F��Yh4R�B����/��9�l`�:���q��*����'��Qw_mIeǢ,����р,�r�7�+�y�b�V�F&}o ���MNb���3�K�8j�����z����| �K8&��:1��S{Q�0-�%���5ɉ�2~M��1�4�,�͖fG,j^�ݒ�0t�g��t~����ІGQ�!�M�p��˕�J�詤��� ާpK�sr�n=���U-!fۓ<�2M��p��8��W �ے���ԏb� ��B����w��&��Ӕ�Hr"��T5�Z`Yv�eg��B�6�^����A����{sL����U�;��u�mW5q�4����J���z�B �2Ӹ�s��	�%!{��h���ФS�bsE�T�i�`�e��9�z1nr�Xj�>��)7�z���r�2f�e^7�$��re?�w3FH������6!ui�%8�G�����I=��:�xweњJɺ�𻋈�c����b�:��jG	�������gofd!ܶЊr����x�7�DՉ����V#�j���pɛ�Q��]��I{iS��˹L���pǴ�
4�:�Ʈ����	�:�'���3�e��˷<{{��Y��#�"��x��fT�G�I�vn�(@��r��qR0��I@JBW�� g[+�$Nw*��'���*l����GB�NE6��mm�#a�$`�E�Z@�U���G/?�!]�K������0�hVqQ,��W�i�w��޼�q͈������9ibb��[f0Sx��Q��IQ��ɔ�~�ۈ�5�`�Ce|����/	U6����愼��Ĕ���V��P����W����@<�>	�_�7�� �9��]�<󷒧�j��F2��v�N9�����Iz߳m�eT�(gHIu�q�b0�ޔV�Kje����j
;?ܣ��&�^H�8;��j��01�LL��PǏ-��!1��Pҙ��&�,S�!vôh��vv�7;����@W��{�����D��~i��j,M=�D-�8�=�յ�F�Eg�F�� r�`$q	iY�\�|Ǭ|�++�(�Jr��s�D?��[��>2�] �Ow�b�.,K� ��00T�����8���-w1Y�Q$���`A��j
#�Ր��r��Ģ�T�����G1�r��;���<�Y�fl� �*�>Y�.Z|TXh���ws̻)���&J�L �OD�Df��� ��ͳ:ڽ,�@U�F�o�Ja��g�į�'GޠC5����)����1�nm���	�B&�3�ԤpF��A-@Fy�����O���(�ܲ�5gOӛ�W×�m��x.J�Gu^���O�E!9�vlӜR�y��E!Iց�m~��;��9R�0`�@ЎF����J7ª?s��1{�V_d�c�u�F�&�+֞�n�X�W�ޏ$/_���8 n��i3ʴ���_F)�\b��a`�8,dEjsT2Ӳd^��2����؃j�F�.	DQ�Sl�_Y��s�E�SH�p(_t�^ݘ��K�a{?$���BY-_` F�m=��Qm̗O�����[�ʫL��i+�3[n�����@�"A�oв���ĥ�������������X���伴Q*'t��a?|/iMb���%C��jk#�GQ욥]BRxHq�	��K����O��'f�OQ*z�����z}��F�Z�m��E`��.��[ם'=��y�0��3��Ī�;, �ˇĔ�0t"8��z:��x�c��>^����,q4�I|�ź�5����%�e��s<h����Uѵ$�3����Z���d7l��c(�(9Aڳ��kÅ=%����@��[��b�cݡ�c�Q�IOj�z�D^��KT��L�����#ҁV�������F��3� ]��q##�E�x	a�b��EY��er&M���nA�k5�bP�c�%��u4�Ԣ5XtC���d-[�vw����C5-��$��MuT!��S�yY�/�q�̄b��Q0t6��TΝپ���t�qY���:�ef.��F8P�}���'�h��|n�*gϱ��
,�`��&��&��?�/'<6�,��[@���ۏ��mO�Q��YJb �_��]/�"�sf�^�/wJ�s'*ݬc�:�h�e�L��ҳ���t壶���滄
��%Y�8_$3�?K���Z^�:��-9	:�I<��2���?��"�T/��J��,:����Ewҍi����i��3�O�v3!�]�f�^���9���c�S��eF�_��*�|l�GS��[Q��=#D�!7�'��}Nv<:'�pW��aǂK��a=x�*����+ F�et��Zd��׸��eT�u���`׸���X@:��6#��U�g> ��Kߧ��u~�>�%v���ա2�=����A���f�__�r ��Ye	'��#b��t�!�2s]��m��R
ǣY��R��#&�����}
���$���Z�p!���������H�L�bhh�1���7��h�:v�0��>��d#S=����x:�֌ ʏGI��M���E<5D\�m�"ݾ1����P��q\�Y2�d;\Vj����!X���H<k��)`Z$j��b�?.��[�`G�0��z�q�x�U�#�8r�F(]mN�(G�-ArB,���k����D�㸟8%x�X��M��q�gP��BMW*�m�S�P�X�Y~���������؅�2�/���ض���lL@a�Ӕ ��'@���1��|a�W�7ݬ�32TdH��D%��7��+�[t�
3w�$�տ��]|�cU�)��*�b�n��
�'�k̦��BqE��0 ?f��c_��J��	��쌲tSB/��E�H.V���	����#�?+��`���؈��wE�G�[t]o@���y��,����	i<Jy�:�_G:����I���t�m͋��SfH�LU|�ө����qQ�
�����Go6A"u��1:�j�у���'
(b���0�7���e�H��"��T�����M�]ዸ�ΰ�.&��:7��H �n��ȗ��0�S�{�Z�`����$ӄ��~���+|2݁��A�����Sd�������B8�5��g �����yZu�a��?�<Ka�J$�o$Xg/#ȳ��Jڠ���8?�� 	�#M�%��׏���ŭR�5��M�u���M[��O<����X>����;�����ߪ�sA���lcY�7@N��"B�4��= oV�HF�`��,�n�N�Z�{��B_�Y�/ �R���.x�m��6zٽ	R�I�@�$ۈ��G��7�W�n��te���6��S?ڌ�~X�u��<8/�K4&t ��Y+��r���MWc�4�8��*���S2%I�p�ﺅ�^��
%F�T���̻?:^�[@�A"�(��&�[iCs.�F�~�*k�p��{Q����.*�d>d�%���}7�|Y3'�s�\�$�z|� ��uIY���c��Vut����b/j:P��u�%81�@����Vq����nM�Kz{O3��@�N!,��缐LWý��3�nwg��F��N&k�fCL���-ƨZi#�Ž׈2�i���{(�-��v��n�\�q�c1���'�э}?�}�M�)��lrH�Ֆ�a��*7^��T	6l+��Ho�E��m��/�w�mz�'�֖�A2���+�EӀ]����Ȉ��ȉ/٨�M���t?N-�6V�4�3`_B���8w%z��p�M\i�8�m���@��|޹q�0V�`� j�g�u�����$�ёz�%��υJ[Si��-A�^Q���Z��G�ɢ��?(������s�8yS���P���g��=�p7<=d+m��<�H�e~��iۖg�����}C�!�K�UF���v�V&:�hZ��?Y�
?u�������jB3G&��c<u��0�n*Sd�̄�
�ȩ{�����\��a�%���S�)��x��(۔lko�x�6�^���!	C*U'q-�1+�JuJ��ǒ��נ�RVd�a�(�˻�y{���J1&sb�JHx�Rc������$V'1䁠&^��ͧ/��v+�CW��Y��rN�0��B� �`� �7�S�W�*]�yǇ��ƍJ��,̦M*�jpƨ����jrM<E����~�>�����00���,�m���b�\�����C�3��OZ�F�)�#�������gO���8-4Dz,�I�f�$JR�?�����Fiq%<\�w�{��	h�	�i��|�z�y!�&��Wѻ}muǻd&	廡/�u������N����v��G�>}K���-�;]A�(F���ԍ%D]�@<A���Qʛ�g�2�c3�k��GF�rov��;���G���~��9��Nem�����.ۥ%�ZX�bV�r%a�˱���5čE���7����Eϒa�g�k�8O��L�Ƌ���K���l�󴭆fn�Ou\��J�ĦGN�1�ʪE���4������6l�(!E��s(�J��A,��ٛv/*"nȍ�W���z�W2��
Ã����3ع*�f�������͔ކqp�L#��\�h�!�tѿ�����]*X�j�F�
|G5�����7:�-�� id���H��������r�k�B�-��m׾?8��,�8��Ҁ�e���;M�e<�v��)}Cn
����Ɂ��0��H �����oj�ȏ�jE���jq�E%�o��h6��Ƃ�s��$����fAW2��X�J���ž��ݶ���	|
��f��^�9֑�tͻ����G�R��	�Xg�q[Ͽ��E^�3�`V+������/�/�\giM�N�ʩ���`�֑�L��K	�X���֎���k܊w�.�O��$��+���r2�8�aYS�Ʉ����:%)3��0<-Q� ��7c�6������QW:瘣������X�2����:E���	�_�����%zjm�=&ےO�7>R��=���m�%��P��w
k&q��U�뼺�Gmy���ݨ�=�p�;_����������*L9�b�Z�?�zj�e5�rI*�G/�C1.�T�&��s���f�����;V�o�+�>de�-���!���=�>t��m����T���i��Q	���&
Q��\ڮ��R���E�	�w�0j�L�7�q�9��v���D�P.T��q�v1SN�?��F@e��f
¦e�Rթ��p"���aP����6�DQ:��v���]�Z�T�r�c��U+pAh��H�L�p�w0���)?�	�:�l�&Ou4Ѓ����yl��tx��u:�kG��"0�ڢ����� �K��|z�@���h�B�x���?�����2ڄ���9ħ
�����k[I=�?V$�EC�8�̮���G`\΋�T��2ş�5m�����w������.B��L;�����9��~�j�
�-y�,z���I7tJZ����Sv�%��z�q���lu(X�U�\X�"�[�?��ߪ+K�]Tb�8b:���^��-�ꝿM��2[�^�GJ$�c�����V�)~{b��Л�S�O�R�c�v/V%�I���AV@n�ws�h�[�/'�S5d*�a�z+F$��y�~���E��ͥ�1?o��������6A����g�v<(!E&��|��RY��}����L�����������:�MrWU2BXZ�	�j1NH�_��q�l�X-����=�w��S�x���A�1a��V���P��
�̭af�xXР����������e�6 ƺ�K����.�2OOU��5�X�%ǟ�3��(ۨ~�g��*&�
Jc0i��Ew�7��[�OBvp��E�O��3��;t�i2��U�X�
����_��[I|�]/Zjҟ1�$�]wj  �5�7.n$m=�@ǣ�MX���i��.2���{��,}ɣ��J9�?� e�3\�t���6C��/�e�a�	g1�V�d삠����_>K~����f���/���Y3�mF0W��+6�Go��m1^��8W-�%�G�hue���?$��Y����A馞� $��J�vW���Zc7���E��ޅ_����^�!��t5W��ϻ�0�9�-J" hi��Pe��X��S��0P�
�g
��z�@SM�f�]ÃG� �U�\iPF� ����P�'�oE^u��٬��N����D�O��p�z�ŝ�{�k{A�+l��8���:��I�i \�j{Z�~�ZN�g�\;p	�[��� ��Y$���z��&���C9���OJu�F��^\�H�� �w��2V��b�rsg�&���F��|L�k�osT�q�����������|c�*�gj��K�@-��\$�oIוV"�x���8�	�@��8N|��C`����
���C�d�����U^�Җ^ف��dO\-E�C����-V.S3X,1����?��kYaJOж�eP0�(�`&���/�@��P�b$=�GM�:���û���iǕr�@S�~^�#����ѳn�9��'����K��m����$(gg5��;?�[X�v�/\�X;���.�Ç�PɌq�Hɽ=����"�FW	���*�}����̞���u;N*�I��Z�e��vU[�}/��zƕ;�����{	���*����>��.e�B����'Ϗ������Lū&U{�7}I;ed��I1|Uɖ,B�����W����',G�[��`'�3:�F�Pj�@0��[<�4�����T�݊(5/N�|��s �_1���Nw̲��\E�hѴi�lU<����q�}~�^��]��켏ӕ�!�Deɘ��Όg �OU���v*�=�'*�,.XO��c�i�F�7�
�:R�aw�Sa�� ��ҡ����
��ja�
U��6��㤛��k��|�X� �k�n��4�>Dv?_���<,�U���+��q���')vk"�+�}s�eά_���P0lXWif�y�9��2�ד~�`�j{G����t��)�׷Z 8 ���I�38-���i�2��i{U�����28���p���-�b?I�AC�&F��ԣ� $�meѳܮ0qdq������Vew$N��#��l�Rh�1ԑ|(	S��ή�!�c쑫�,ć_�&wY�*<��4�I!ǎpOkl����p�˄�/X��
��b_0��AWտ[1
�j��ef�$ �5H��P͜XԮ^꛴
���@�]G�ݙX�����C[����l������I���v�/o����h�6���	Wd�n֨uh�2�D�
�|)f�� �#�5i5�C�cH�rX	�S0ȭ	 �m;r	Z�O �����N�Z�N5�5���.��}F�˱Ci*���,ne�A#�mݣ�c�-�x�|�a'U9۬)��w��̥N�ڨ /�_ �]��_ig�*�
Nc���Q#Qe��Rٿŗͪ����k�gA�1�����Rb����0�y�/V�Př�(��-���o)��ɏd��pgZ&���([��F�F<.W9��n�h���3H��i��ˁ�a>v�5�N&���ܞ�HR=0�e������@ȱ=u�i���Fv<�\�gXKG
�7��8�V8��7�f�ݜI�!�2� 0��ם�u���J�6-��8��哂�VW���]P
�[o��A�s参E���X��
�ؗձ��^�N�P"��eel?�k�9������@]�>P�W��Z����N$<Z��>-ވ
�P�]���4���U�1 \��
pcbɼ ������QmPʬ����.���l���pz�t}�e�"��c���P�8���\���&)��s������ڥ^ �L�Lެ����!L��8�g/��Q�@R�I��N��I�Ѡ�y�JDIT�ڠ�w�-v��V�Zەw��ii�E����Η�)��7�E�FFK��D�_N��p��#@'ӁD��ޚdE�N�++�{��y���i}i�?bҶ����/���� �����	�@�q�,���v%z���]�bʜև^��V��j�_C���e�NH�ը��+1�[ .o�!���E���G\rX�KmJ�j& Z}u��M���5�$/D�� 8�c�!��w �@��W{����u���l����#B���֕m�"?�H��5_�
9ch�R�xt?Oi�Gș@p7Ɲa�D��N�H�q9,�s���z=j� ����4��l	�����pr��
8�c�E�;���t���[�w��kMm-�K�m��k�2x���.�e�Z�����SQ�/���0F̾�����g�����ag(3i��	�������=`2p�­�}���8�u���y@⒲U}�[�/a~/�P�.~��^S�kS~�M�|�=jM�\|�遹���;!#:'M}�u�>�"�fpMO.L(ۋܡ��B{�A �ZɕbGQ���i����^�S���蜼���R�/T��M���a���:���Q+	|�6�J�X"'������82i�~����TR�q��?�r�����K���MW�����e���ѡ�N&W��.j~a���J�a!>�o����ǽ�+u����,�q{vn���F��ϳ��ưl��41�Ԇ�~�]g_J���1�2�w`�q{�kP���ⓐ~�o����K��a��Q�]L�B�u^����`+e� �Vl��\P��8��}N+�@��U�0A��	�#Lk�vc�\13V��KE�B=���@�P�E|r�%�d:V�H��tVO`1�Ѫ��
3I��Q�D�F�IBؑ�&��p�j���Ue��-�/]�U�D��Fe@���kz� 1�!tvv��Wj�mWRo{���K6�FN�n��e�-�f,�W�&E=�t:��@C�&'���]h>/����C��Ӆ'p5'>�s ǼTM����n8t���$n���p�&o�N���2�1}�K}+a�O��������䜩�aRd�([��1�|�e��g���Q�N"��k�7?2O��j;mH��>��ү�,����fĭ�|^G\}MZ������o�ULl���z^Y{��|��� ��C-v |���a�4��	 !���f-����v��pV �9�h0�?�@RI�Y�M��F�9��c�\�+�B�w�-�^����&0J�2��O��tS����Rn��q���9$�0�	��W�sX�Z"�����E9��I}A�'.�N��gj�'�����p�d"s��LK��?	r�F�EO������8/��җ�5-�R4^b(�G)N��ʃ񗶭b���g
i}�B�o/d��V�"��{�!_*V�曠�������1[����d�(�/���,���R�����k���Yg�6p��OdVR
5�j��Ę��:�Ŏ��Q�:����ə��
aJ��Z�l�9K������Fz5��h �ZCv~�zg	��Ǌ6���T������Ll�p�T�<ͳ�����@zb�N7"���|�p� ��.�Vi��ZRb'��<��0�!R�
�.>BqZ��Ǐ����P��z����ƒ��e�����S��{WE���9��>[]���%��O�XGr�@r���Q���V)g₥B�Snx��w�<9��Jd3��HmZ����oΉ��8ۘ�5������Z���=�+���do��L3-���e	�y�ǔ��ۿ��i��@)ܪꏏ���ˍ_T�ZS��
�z�3�ұ�
?f��Ǎ��kR<)k?|��U~�}����#�^�{�*�v���y<����ð@��.�G�X���,m�v��a9/����@VeN'�c�� �Bbg�*Ͳ%�&������:W�Q��S	
�S�RQ��A���}�'�v
R���!��u�D�9��B�
_�}�4P�mI��E����_�����8K�'	y&ĆB��u2���.�� I��<9�����d^�dSi�j��],���}#���"��9޹�(ڛ�P(��ề�����TK͖l���?���p\_�ti!=��V76�Y"m.�9Rv�T˲N�X���q]a�Dm��c䢜|%<\��uo^��+w����"�J��XN�R�>�� N3ߘ����]�I��߶A�����!q��B�}��׊Q��!&���Ƅ`�����C�N�ll�'-C7�楀L����ĕth���j�k��=�aƛ��� s��Q�#2 �Y��¡�B����h�VZN+yL�J��N��'���k��9h�m�z]�S$��A����<�o�A�"��f��5au�.`�2U{�T�k�^� ��i6����Ür�;c�6���9��n/�3ѷ���� �U���b�Y�E9�HM���B5��6S}W���'��cϜ���)��.��0�����6���Ǆ'\r�L2W��aw^��RP���ְ�{�K?�lş�8�+�xv���I�Dax��og{��O���&��H7�! �ߗԞZ��,��IӏLő��B��c�����w�W` cJ ��ȩ ��y����bƔd���o&X�!��R��KЪ�!�AY��uk3Lk0��X�q��� �����$!�5R8�d���Z�U
��Zo���a}.s�����f�g7%N�	�q&GrP84@O��z�f��Fj�'���G{���򐶸��@ƫ�j�<'��T�+����e���ΐgQV�V�j8��Z����>k)# �m�^��CP�+q����~gJQVy�5f~�?��[���o2�)lt{���rnIN�mɑ��6G3|v��">�7Zoy���O2�B��%�5F�>+u'�J��H��=�6>�x;\NSD���@0�,$�"�����=_��E��*�L口��B��s�G"~o8����P�uz���7 ��|��Y��:���O���Y���H���;Ŗ���1E��r@6p��<��n�1dvh�g��V�ɱ#s�Į(����}M��Hz�-���|��PhV��`�*�qa\5����-7��;9�#��Q��	הk�4$�Q=|Zì!f��]��MU˅�3o�z9�"Ŝ악�A��:��ԓ,��$��3X�|!ѳ[y
dmY���Ǳ��Zu�䀽K�L�U3�Y���*O�}'�tS�ן���x�(�4~h���m�<l��}����N�I�&*���+�z���SL���F�>�~=ǀ��=�/.텢�����TthsBu?L�I���^-!Ee.��?���,e��5���m�x���1E�;SX�ɍ�����-f�N!aT����x�E���%E��+*�;NX���%�[�N����mi&�A�ta���@YY���Y�؊J
�� J�]!��+U6nǷ�[	�M��isCE?:[�i�s�o�t#OY�.e�Ea�p�4�V����K�&��r骮a\q[M�k����sY��7�����X����d�W�IDd��H�S��]����XI@_Bv��@���i�T�K´:�e7G�V��A�i�M	Lvz���aHn���cA���I3�j�k�%��Lڕ�/CD�|�������@�d��EX�ґ���,���h�(�7� �H� L֓��B�(5�[iLq�ڿQv=ߠ����f�����-��DC�P ���=*����[��d���g�K�{Ó5߉?[?��BE4�]|�����U$pxI���mM봥�u���NˏZ=�f�*I<kPoU�]LoB*�`�5/ˉfWy ��8�&��C�Ҁ�/es@�j+�A��S��;����1�C�s>���0o����Ɠ�D"��4	��Y���GNv��T��n`��~H}��Cb7�c�V:�7����]������s�A������'���[<<i�5����/0�כ�E�U+'1��ڧ����`y��P-�����B������O]�����_ M`cv�T���N�"����
^ؤ������Q&��ӝ�"Ԁ�rT,!�ϐ�%"�8���'�	\
�-�[�$hzUf�MG�$��#о���V �$\�Q�MK�8�Ik��-�gQ'^�w�5��/��ſP�JFO��
F	r����\�[�^���֭~�����*wLbl���ʰ������Xg�&��Ɠ�{�J���6���,��_��7�������gQS:���y�3jU��ݐ.�zvN�ەi=R!nc@��W��(��z�/*)E���H�
����"��G4V��;�]u��r�p.��b��|�6
S5�m��a*��n�*Yxej���U=�}�*A�IL�d�����/���:��좭?�jM@�	�}6'TD҅�˃�an���͞d`i�23��-�%XK�B�aWA��T�⊕�jUH���;C�+`G_Ad������i�"Dq�gArE�7��HY9�Ñ��جA&e{"�A�98���fY'����7|�^I�Bj�M�Aw�T���m:�j\a7��>�]�#w^��g"�@��Q}�B�xd`$��Lj��$������x-�\	���>���c��칬Y�J~|�Y�����S��?��5����=��O3I����a�?��T���\�����=&%�|�7y�����k�re�W�Hx�5�r��/�:��iW�Ow�WZv�%���?��C0�y��5t~�\�ǽ���ַG�gz��� ��ǟz-�Z`�G '��_ �v�R������6j����O�*���dR/a��Kc����p	P�:f�x�w�P8ǽ5�x�Iw5n���~�V����_уtM�ͩ�'�5�u�A\FJH��\:�7Slǹ�fT3lHS1�
��^ >�V�g!F'1�^]�Wy<�o,�)�G��_>4 �ލ�u>��I �X���D��S,���1UjX>ۊ�S򶘄�|ue�y�i-�Fk�JSS�w�����L0~R��ٟ��B��Q3���Г��/ ��n$�oJ�{����TeB5A��̆a�Ҹ4�͟����:�=�k�d~L���z��FP�z�m�b��{tڝ�TP�G���]�I�A���Q'��O�3x���jD��é�%`!�\鈧߈��@�/��S#�@2�oON�'��Q1$�w\�R�m���L!�}z�H�DC�1
�R	�-���K���A��(�g�(�� w�e�`F�ǿ@��y�U�Y2��$-�G�%[1���X���4(Y,,_I$��=u�җ����!k���e�^y`0��5��i��4]#�o*"b=�D�v��<�E��E�Vr���:���'J�k���)�J�I	�1�~�AV���lm6�zת�,�V8H�0o�m�t}�G�Y4�v����O��:|]�[���[�n-�:�o�/���lER�**FXn"���<ֺ���~/�`��j�ē��Q*�1,<��η ��H�h�N�sp�<�-�:�u�?�u\Uי�i�ښ�Hq��hg�ů���#��Bd�*(�x��9C��Ӧ�, u�F��k����B��ޱ0�]V^Dzr�\�>����[A5G��D��Ȃ�+E�~�ɓ�(:bAs:�i*z4�PJV%QZc�g�J4icH����Z�|hW�X	�F�4Ϭ���/�?n�m�Y����|MO�_q�.�ir�"�2N���|J:�&v>1JG|�
���r=������Ɗ�b�Ӓ�Q$�mąt��<��۫�Ǒ��Wt���:b�KS 5fH�y�T8��}'�'�|dL8ᇾ��trr���1��#��3zl�6�r��U�XK� =�i��� !�S�s<u��0��k7d�Ӎ\h�L䉁�E�b�x==�|'�֕6H��Ϲ�d6]�h��22�Yţpe5�b��p��9�y@X����R�E�p2�_�B�L�VjZ9&
�8m�nZq�f�-��	�8�V�g4�Y1���sJ����O_�䒌��N�ג���"�@��}�{�/c��Sd�����C�T]óM��W�o,�7cd���z�nlqblɱ�$�tM��#0����Eb�Q�[�%��i��_5�A�i��q�w�<�"�h��ꄧ�zd3��X!Rk Cm݄k`p9;�����Ԙ]��z�[X�kp/)Wd]��|���}�J��p�TA�W��@vM7�o�ڎ8J���������mH�o�)�^��Q9LK'-m���+&5[��iE�&��'��\�	�� �r}竝�q[)����݃�׃�/��Ñ[XO٥�#������^�,�Z6D�
��㵗��2�0�_�1��Gi����l�<�g�R�x	v��Z#C��W#��I�Q��N0�8b���fJ鄠U���v��;��ѷ+����r�A�<���Լ6>�Y���tq3nl�#{�T!�������!/���B���ͣ:<��Ka������-�0�G�w ��t�n��z`�q f�5�]A���.�0}�3� RC%�k�_r�f�OVMN��V��2��.M��T��Q�z��[w��Yf9�)����@�E�H�ز�)RҩR��U��/�@�
(�"ϒ���`���F�*Y~wdv#SQ2R���[2�7�E��� 5���8ɑ���Fi����}��;�x\�Y9	��s�D��)���@�Bpi�c83ͬMy���I�3/�ς{�M:�H�RQt����X�����;;ˣpQ��hfc���vu�~����� ���t�cb@�*�4+l̂�jk����w#�2k�S�K�rJ�HDs��0�$x�x7�_t�4���Tx�$�E$>�))X;�)!�qO��Â�%,f���awi�`KU�)d����L�=Ѕ��	}�Ǔ,R��o�QC+��E<�an�1`���^�ɸO�	k	��}���>V�M�k������X�Q��2���3(����hO��Q3iY�,1���E��3�Y����u扁3��`� �Z��`/��d����NɵAc�L�hE����E�������򠧊����_�#��KQ@:�L�r!2��J��X����(�wB�ު�ouj&�C�ON�m� v���\��c�]]��:�ଜ�G)�@2m���yGV��A�k��T]ŁyHd���v\�O��5̝������~9�U�v����ny"��i֊�G��ʌ��~y�5�H7�7i
[�5}�u�d�����Dɹ��9�-�'фqf~]xP��Mʱ&���t���j7��_G!�
?�bOqBe���+i�J��~X)�mt���ߜ춗l�{*gB	��^q%!��pd��8-����j�;��9Vs��ׅwOo|�x�:wI@�S�ҋiE�,�b�*� ���7!i���X�]�&m%-�P��*�o5�`��>~�$!Hk��R�bUt Ԩa;�U��+����Q(����3���t�a�F?g� ��m���V����R.�6����m�\.�cyX�'G�J�>�1���py��D�- �u����Ԁ�B��������Ho�Sz��-�/�KK�{:crq��:z	{75�Ř>`(��������,@���	���'��6���r9�\W�i�Wu�/�y���e��B K8_g�K��k�]$f��wY�h�Z�PJ��~ss�B�3��?>z)�C���yk�
��w޳*�E(.'������ !�I���� +�|���[Z����ڙ�{��w��C��cSM��e�`�-ũ��h[H�=���Ȓj�3�)�l�b:�@ǽ�o�}	�VU���팠�E[h���p�2�9�?�����˶~)��0��~��oM�<��V�]��+��@BYZ!C��`���|/��I�eA�`_�T{/i1w�\��UNAм�n��v�Ib�h2(�\�p�6sy��H"�AѶ�B�fj�0�����S�j�n�{?4�\��t���M@�B��hl��"j�>rЩ����j/�˲q�Z�渽�}��Į.��-g'�f�O1�y���9��/�~���i:��Z?ȡ�+����2�q�ca��j�~�l%a�^>}ĥa��$�(�ot�N� !��ay��EH~����𞰥�8����p�������^���,�:�DC�]̦�@���¼1��J���*^�K�ݾ�=i!�p��߁���"(8������e:����b��w��1i�M�.�$��)'��5�I���������%ڎl��++���d�y��'�?j6�Bn��̌|OB���������T�>6� ��^`�_���b%�o�T����E>P\�f��u�"��c�y��H�L�!b�l����2�RL�:s���6�b �7�F��C���Ad�i(�l��ճ9Kj��ߔ�X�V�z�Yu._s(e�p_���0+�H�d�i����ߘ������0�e�%�jꄿ�����׹�m�ܽ��z�|��7]�d.� y��D�9n�!���p�D���O�G׼�a/����?�N\i�)�����c�ʥ$�y�K���)B> 9�@��_^ϕ�sN>����ߓ��V���Na�9"�qԌ�+�y�!wb�b�h�5��@V9��U��� ����ڤ�	����~`��o���<N	t�bDۑ�o	X����8�oTҗ����h0Z�g��攓=>e6�U�\,`�(\V��ݟ��b�&����'�LU& n4�� qE=�c�(O�P���s��X�QI!�h���nh.gC�4C��/�&�O6Z.Mr@�[��	&n��Y���S �V�j���q�����!��˧��n���>1�b�~4P���C�M�g��V����FdJC�h���z�(6�_�
�g��$�(^/R�L*�{�Lc��8�V��2��^hf�\��@�7���y�c<��f�e�y}ˌQl�$��VM$���B�/F�`�����/��HA�v��2�efS�6�01�s`�lQ������kq��Z��{�Y�z�h�9f�޽`C�m�����d��*.{�	UC$L�-&�E?P��,k�еe�*�R�a��ѱ4t���bu�c��.w�'<��h�z}�8>�=��e`�<8v���ېpy_@~VF��4	�Sz��jخ� ���kKtLK�!0D�n$��Dt�5^2�SW��ȼ|�	@G���P.J��I>K��0"���o`�/&��~5�hv#8�4���C�N��o����8[���ȗ	r�GgIR�����U�-�F��6��i�ǜe�)͂㗘d�W��
Z�W��iҦ܇K�z��P��Bh��ҜQ�Զ8炎�[���0����`G�8ʱ3�m8$�i���̌��g9�ˢ�׳.�_׉̏�U�S�:ߧsX���K��)!L(��4�{V���8�(m�Q�����q���5_�^
�L��/7`$G˕����+��}�x���`^a]�_��"T�˸����%�<$�} g��������D��^d��p2��7���:2�yM�
��)Fj��<d!��mʤ�8$"[j'����	�je�-����K��އ?���#0`�vC�DX���&��<����A�z��֓������d�(��m�*�r�R�Y����8"? uY��$D��^/e��)�Ґ�� z�/�%����9To��cf��
���u��ק�a�����TC,	�!OY&�J�Z�#���p�}�@qTm�"c^� �~��l���Ҝ�O!�9ܞ}����z��M\c�f�#�j�G��)hnփ���Ő  ��&��}JW� ��(2Z"�o7�b���,���X���`�d�bWБ+�|"��Hl�7֩<��\D��6���p��p#qW�v�5�N�e�s���m\��RI�
����+��H&�-�������~X�u\��J��*�1���mSO�����E�0l�	_-c�	�5^⤲5R؛:<�Eb��n��u��2ty]'�����4��?�$��Ϲ�{�����n��/�����{�J��$7�k��1	�lE���Vߪ�.lO�{�\2T)� 6��3�L�#��� h�S�T���ks�$ �p�bU���KT�i��J�l���q�|@�}XL��\�N��/�x=`�$e��ԫ�Z�Ur�z~�fs������t8:w�z�n �t�#�0lp�V{֊T�$~@3N4
��������g�c@��TQ�Crc���8�5}{;tv�E��	.��N�]���s�E��3X�rV��?w��+���!	�����g�j��;^�:������03���|ݑ	{�w�1!n�z|��j"k?��t_����.��5��[a}�`���9���g/{G9]�1�7c9��
e}p�
V� �@k[�^Q9�<���7�x�&��^8������އ�`X[��4]:�X0J^��8V���ԙQd�m=Jf����uC�� �%�� �ߗ55�p�ENml&�'�oq��:~�	!�OF �Z\�}�׃�Pfy�s����jZ\+1���]�1	$�<�@��Ѡ�BFli�4��l���Gj��"~]Ns"+�h��%+�Ü7u��
�A�I��)P��΃��0u�˄�3N��
�lCU֝����}��  	l�Ge�9M���J��ڍ�I<JT���L��s	ax�jKΛz:�M.jlR�i�YhK�5��Z<���|���s<��H�9�4��;:1��q? �
�s���+R�E[nuc�ۋ��rx� d�G��am�M>���؄#\㾾�<��kOW�(���.tE��0^w-�t��
O���<-i���XSF���������H���8	sl�wsʡ�U���{s�2��̕�$n �uO�j7Z�w2�j���EX\q���O��(�v��ꬵ׏2��%��L��B���nб@?���1G�n��G�]�=��)���{���d�*\W%YG|�P��O̢�#�8�!!~�d�������/�b��wd�P~�:������I���`{�����+jRlU��視~�%��l�T��tߐ�ݼ�Tyj�%K�>����t����+�v��E��>�6���n�Vy�U@Nc]�Y�!�s�ˉ�r�|����ͮ*
�i�`�6�m	�1f��� �B�BY��k�j%����X��M�{-�"l�/�-	& |��ʶ�ax����!&�d��$9��?s��h���z������̛��X�7�Ao�`�>~֊a�mJH2,��>Z�pX}1zvFk$�v�@q ��t�����R���y}���V�����N]���,2|2���]Y����� �ٮH��IC�����[ɍ+��?	��Μ�=���wNF�/f�s�����ϞR�ڬ�[��P/�N1T�_�a:�G����Qᨙ6����(\�{������΃H����4��ÛX�o�T��r��c��//!ZKZS��Ș�:���޵��$ȱw7�,��J��). ��5[sS��kPas�(6���p2���]^�s�D1E�H-/{��뮫|)A}����/hX�?����r�"%Qfg���"��f��/�ϙ�����f.~/�1�~����P��`�H8˃�y�k�i(>ޗݓ%��{�}(�2Թ���y���)�M�.��\��x�U2�h�rD~�'�^�4�1�y����v�[E�)��6A��Ի���Dc
Ϟ 	n�կl��e��;?���+W�VZU�:y?�v���D��5ԏ�,g��3���ӿ��<c;��[M� ��W��b_�¼�;"A�N�;�.�cAgk/���SIMu��!��{=���JYP�؏��O�~w�Yj��5�r�˨$.Ѩ q�BP��M�j��dK���mx�����!�rL����V&��7Gb�Է��zr�*�?��%�l</~�c"��g%�����tB����e}��ۼ��B`<���l�D��f�!��l z���z[�Ak�e�Z�D&�/S�q"{�q}7<���De�:b�Zl�"1�� ���U�F�i���
�v%���$nAF(Y%~���k��򔛐*�\��յO�

øR�B$���&vP�]��������c��'0�0�"hx��xnfЯ]�X2m���;����fv�D�f�}&R����f8��#�eo����;�O]$��A�� /�7I�
����׹:/]��b2e�@���	�k�\�d��l0q f���wC����~_}�>\����	��iy[���m���ҝA/#Ʌ_�~����Ǻ�0���@fB��J��0����T��̮j4\��_��xҍmE�1�m��G�'e�3�˼0+�{�Fg' I��E@�7��g|�;(�`�\N���RW���R@k��'X便te�
��9U���]�B�q��ti���LD���
l�F��C_�����H��T��Pm[P���~��8�T^�P9/��m�.S�R� ����A���o�NT�iv��ܾ��Pn�Y�n2�J>Żg$�'�a��
ʥ}��wM�0*�S<�Z<I+����;p�.��r�k1z��I���~���9Ǳ��m^�-�Ĭ��W�д�������t�Ne� ��o)^��(V�@��i��[V�jA0yX>l�t|�l��tƟ[u��]|�V*��`غ�r�1��#�*��[̫#h)�� ����V�������fxą� �{�v�"5HO�Cm+AaH6���~R�8c����L�h6cp��!�RP��6�D7bז����3���K�:�� �H�>{�:{Y��_^Kzb�F,w6�*+ԗ�V��ŵ���"��j�.� �+�����A��cqM�q�\��F��x�lE;�d�6vo����y<7��������h�8�7=��+1�勑�'���I
X�e��^6�9�$��������� "��,�:�������G��Mf~�p�(���lL�3 Ќ��A�T �6Dw���#�9Vm�y�A9l�΅}Z;���{�	�����ղ��Q;�<^ˮ�\���-"�Oq��͋�����&s��Lf!����{2��A1��C!u��c<�G�b(�r��]��ߓ�N̹:ވz?�5�r%�ҡ�Fk^�����3C>�X�vw<�U}q����mۆ�vd�Y��r2��8������a؉*"٩j�X���r�Q�-4%G��öQ����U��_���6�b.��A�x�]9��&�c/�I�)Io�J%g�� 	�k��Է�_�<��ʙ��&~'6��W=9�mj'v����`�8�xA��xg�\��B��W9;r���|�֪����Q���\�c!�J5V|;��Z�@���A��_J��%�G1lSj��{QI�nP�H^V�HA�8�ء+�&�8�c���&4w��V!��<f��y��P�����R.X:=.��v+�|��FR��*��Ad���PX=����J��+N@�2�c�Rl�1���w�x�$���?�TH���h�?��3���.�V�,(L�*��" �p�2�?(L���h}4?�6�1nJ@.�/]��¡�388Ǿ��ܥ�R���d�f����Q�v��oi6'�AL�8�oCc�)�H+�6� ��R�p�%��!�Чx�K�������;a�ѱk�2u5r�����S����_΂��x���/<�|�-$:Y�J�Y�m��-F�DN�'*����Я���E2Oy�O�9"?)زɊ�ެ�s��%��t T`[f��x��J0�����I�������	���X���X4�����G�f�q�B�����CH5D|M:�Z���RY�iK�.o��*����3��d�2�ؽ�x!K)h	�F�rc��rNK���w��x���������, ���h��nn��kc67�ӏ�g�Tخ�wr'&@�le,ԡ�O��|���c���_?�s���f�v���)�RmL�%r�p;��o*ƦaUiY5��9�7�����$�n�ޚ/�A�∕/��NP�L��X9N/Q��O�ݚ�[�W��h2�*�Wup&X��i�:�����.�����
��P��v�����6��!q��7:�^O-�<��JZY:ޏ��zKS��C�Fd"�<�r��Yl��N?9;~I��^��n[g��*g�ebK19�9�Z���z�T�FDU���\�"�yyLPG���a�b��wd�5o��c�<�Y����I0�N��(�^�81�������_��D �(��Y������03��
[U�`�p�"�Ο���E�X��As�c4��枝孮�����ꂣnS��|+����L���*�ӭE9�����pCCgg�%�q8��2��(<���L/��6����	K�qjƛOH���T�G%����Fǌ���=�O�I&�Q�IYW��n'�:ѼR��A���6��F���?��A��3/��A���a���$����'c���%rT�����ts������f0����Z���fR��t[��
����_����<���T�t��`|��ʖ����I��$P�D�Wt9�~�(�+��� Nw�k�h�o�VM�聠�	B��?���=�f���uIp�ɝY5w<ZK�UJ�j���,8��2��B�|nU���'1���'�+z<|V��D�>�G2M�]�l@�!{?ˈ,���
�	�ַ'��;-�L��*������\�W~6��j��~��b�>�g^N���\�#i�
�ui�����0_9��L0W>�5�wKhF�f�����7V		1�l;�A���Y�qVV�<�@�[�J�>�?������OY~s�3یǁ𱟠g���B�I� ����{⼓�dX5���*�k��ӕ�(�xś��r��a�jv��aӊ���i)�WF���ע�MfY���ڮ&p�Q�<���6��o�
x
�g�B���K'[�"g�M�G)�f �zt�|N
E���%�Jv��;\�t��.��i�ZP�[����l�
[�h��P_�:�@�z��Z4��`1:��؝�M��fd\<�n�dFL���������5$�0��4i�eӀn�3K���$���WL-���WC��ɢJ=%��[{�h���d�y�d�����O����PZ��lCy�8Fw,��TL�AՊ�K��glܐ?�З'�1<$��SȠe�D�<���1;���3n�⣌�l��b�W�c����΁>��H�_~f��{���9j�Bɍ�W��93�3��+��%id�S����4<òk���]e�2����қ�u�.C:7#e*��c���#%Z�7na�
����j�&�:e��ؼ�""8K������j ��n�������H����D-Ehz�y�D���E�J�P�3��{\�8ͮ��K��F�\\��'-�S���`׉e+��IHGk�ӣ�B"^{
>N��n��!ɰԗ������Kw���]T��rK�xHG�3�Z��.���5��;xe��m�_9G���!�o�Mr��}�{�fi��ƧZ.�U'�4�U���?�bd�H�+���v&�j�>є(�mb�w�B\Y�g���n�C�A����l��%p=��1� )��2@"�?�TV��G�z*�%/�I�GH�[���E5	��x�c���X{�G�b�)|��[��e%*����YI��^��¨��>o����5%���.vF���[�j]�"1Y�b�D4%��w�a}'��Ӣ>���/tu|����ó~_73�7o?q�Ao����#���+$1�b�y=�Xm�<x����$���5.t$���P�r�?�nY��<`$L;�DH���rh�}���JE��8���O
��Ձ�W���q�s��׵#�<臔�𮮏�N��t�mxd�]�<6��H��[�B��YRN���Ek$Ɖ��Ii�*��u�R�G�����L��0��E;�:�v���^�Ga7����){��uJ���?�V���:�.�ܼ'�g,ͭ��E�ٱI���W�M7�t^&�8N�P�ZV����������o]�V-!6�\DX����R�5����,��o����=��B^�Y��a@
R����3�x�'�ocVHI�Tϵ���vm���7��)���'v4�^7����	o]���Cn��[��f�+%��ŔҌ�kw��/KH��mA�����}�Y���ixEO�����́ȕu��ħ��&��އ�ׂ��(�滩)��RZ�~#4���B����ȫ/���1;P���n�Ӛ�jL��4[T*�ݧ��l�*��7����x����G��pUA��X=��^se��b�1-{9��$��$��;I��*Tsĩ��ܳ�[ҽX2�k�3W�9"�qW'��a��yӟMc��b�޺��]��e#��X��x��!����'����Zj6ҽ��"̝~3{�W$i�/����2m�JH/X�4R5��ò�)=��fn��"����<���7�d��;�	��8�u�N��0L�F�ḍVE@MF�I��O���O[���,�.�=W��Y$*`F�+�32tJ\�	qG�꣌�l�(0`И��=\*-���i8�s�Aw"���*�b�^Y��ב��	pK=)�q�C�q�{%7
^�����l)��T� �`�0I?6s�����jܜ�P��T�L�P��r9��U��N'�:��=�61�̚��F����lxϡr&��xF��d 5�g�H�9��ϊ�T�$�u�qsc�]�[�(�6s��L���E8~���+��b�����ڂ.Q� �r��yi=E�!}��Y�*{��up�Z� �$ߟ@��KP1��o~1�Pwq���V(�qޥ]r���>_��?fmj�L���"��b���S�E����/�o��aP3G�������a�+���E�u��*jOݿ*4{d���"��3�i�?�!C%Jft}|���`~
�E5�N)����Lh�g��Z|��UB0jM�����w���:��F�
��K��דP7H%���8�Ii$l�����̬
���?ͮ��$X����uX�(Y�S�j�%�9@I˴9�6AܩPgF��&	���ۓ*��W���+
��WI��#���\�G:�lI��{���Ah.Q����K�[��#=��b�p��L�)E�rt�N�,�d�6	�oIa�\���of������?����R�f��&x6u�X���ԏ����&�稤Ĭ�?�MO&�0��H��b1�oD3��گ���)Kâ�
@*��3dR�mdF�����u���B~A���a���y)"�!"���P���`o8�*�� j��u�����Rzb����K�m���0R�A��6[��������߮�~z��r�T��P�m����1�?������Ѡ�d�AQÇʚ��|IB,ZE�����ʲ$��DbU����@��fM�Dx���2�]j�5܏���!?��"�I�t�i�5u��@��颢F�%OF{ 
X�(���&	^4�l@\�A�0�)¢;Y+g>A�x�f���&��?���C��;Oa>������>a[X�P]O
��%�r����y�O�n9'��;O�igH�n�&y�zĄ(|Q���~܌�I�[����3�����AF��z]�1.��Ԉ�Y��STqa�2
h��vB�aP`���xw}�2��0��ْ�Q_É��
Q�̇)h��Tw��ӵ�?qރ�Ntr�0�=\�tG��i�8̼_G�d�*O'�<�T��D��ɚ����U�� �g��(�gb4!z���ji�4n���;���Ҟ
�����k,�FZe��<Tޛ�R�8�'�CAD��c'���~��{/u��Z�X�X���v�%��`��j�bh��Lʓc�,�㉵��`7<mN��NޘX�(vj�?�NC��\�b+��#��8����A���_n�0����>ttA]5��;�� �O���!_�+�?���>�1H)��v��P�\F�(�ˆ�Tr�Ldl��Mϸ.���53��03���!��F��o��ı��a.����ӡT��dcaT�o�ļ�!�6sw��<0HB׋R��^��W>�ӕsX�~�,u������߰vr���ȁ����|���
A�����	1��O1!�Y���N�������Ih�=6`S[����zw`2I���K���l����w�d��������ܵ'�±�����[~Ph�N� ���Y����\��VVɂ�����{�s��o�-%2��G$�ǳ�
P��NJ\n���942H �g�!?hj[���sOF]/6�2�jF�����|�d�B�qd5�!"�(�x+I�����������oQ�H/���U~h�wT��đ���� &�;���ڳ�z*.��Ŧ>��*�qЇ�v�B�Z4ceA����K��{d�xO��v4�L$���|md!n�|ФULAQ�3O�A��^f�feI�Ѻ��o)Xg�վ�e����mٔ���o{���M��u<�(�;ا��ޙoZ&���B�~SO�����Ƃ
v���Xd{���E�I�r���k z\��aY�}�=�Gu���3��_���=�	�:�A�J�<���wi!w�N�܃x��Ġ#P�[�LN ����p�}�j��{Z���
LH�d
���If�(,�An㢇[	��x4KR+Dx�g�޶є(M"��w��RVP�%�T�⍢��a�>��!j_A����ty�nz�Y {�[k�~Ȣ��N�'	�^��@&�x�	��@��oEH@?��zx����b�᭓&y��P̓�����f	R-��P��nt��Ɛ���`q��NX1Q?�ѷ��f��V� �j��	twL���ǉm��Y��_̾oK]�O��%���|Q�{%��*������r>9u�m�'��|?�ƹ�%�R��?W�0��CeBx=�)�as=���0�s"縟R�\̢�i��'���5���S�P>c�/螯yǔ���]��2Ƞ���"!�sLSl���`�O��A�jh�A[���%m�$��4$f�R]�2�����f��t�ˋ<�rO!'{����"�b���,2J��ė��3����[-L��u^����0���?�����! ,�y곍�ڵ�����1ȉh�����Dz���{�	�/�x$�#���^�I��1��f���ۊ<1Y+{�M'*���)oEp,�ЏeY�2,P��|N:_���~�)-���%���V�r!c�����`hS���I�&��=6� O7�&yV��r�������r�up�l�X.�Pf.1R�	_��>�}#�@�h9"vǚ�C���@�2
~)i#�y�q�	�|����W�Z{��"[���_�d�);6t��n��z���W7�4j���0�)�ð~��&�oGoz7��Ϯ�ǽ��Ym��ƺ<@��C��!�am=�_\6^x	v*|W]�7ؼvT���$��>u��܇Me@�+�=T�	����,(!�k(c�;iC�o�P�{+{�?�$q�݆H90�OS�ܐjt.엎`u��@.�V;�ϣ�f�=JGZpmA��U�De �e��]�_r7�&��su�C��`Fģ\wt���R�|�]:J} x��r��$YEv-W��is�vD�Xrf�9.6�~�(��bR��Չ����l}�(t�Wn���د+K3	������n�y��ؿ�*��<iwѾ�&�6������k���?�]H4�{��.��/߀OIB��k�f��( ����_�gBԸ4��anb	�^����`�C+M�Ѣ�XHw*�#�ܦXs[3k|�>�����v��}�}�f5�5�?��6�>��\Y���E}l�2�2��Mt�@��$c�H00�r�Z�fe�>^]�E|!ȣ����*�p�m�&[o�lPJ�H>䍤���Z��%��(4��h䛊|����|�ۣ�3�)�QNKM� ��v� �7aM �ݔ܇v�/ٞv�ɐMh���42b��%N��.o�U��8����� �7UDÈh�Lϴ�c�_ ��	@�I�	�ܵ��m*�/�cCyST���q�S��\t0�`�:�~U���mκ���ܹӻ hsĜ*�_q	�yo�H�p�P4E�?ˑr���{�.9�6��4�R��4_6�ö�4�h`�y%�Sص�' C�����Y�w������\�cۍ*�"���u����Nǖ�zf�*5A%_�4{�^�i+���tI�o����=�3�o֞'Y�
�E�|-����Đ }#-�`�����������c���Ѳ�ӎ��4>�2(���w R�4IPS�Kmԧ�j�fꛋ���1z0'}��̴2<�[����+iӫ~o��w\��9��A�~�f#�µ�<�_�\��{��s=u�ھ��_"]yۀ���?x�����+<B~�M�c�z��Ɲgw�4h�v��!���{5�`����ì
��uѡ�w��2z]�Nɩ��Vt@h�0�۳p���P$�����/�ߐ5cղ�Z����+-�M��  ��K��%�D�x��&�s��1�#Q�V�~�
\s�ؓ�0�荶Z�4�jew�E!���zvIb�Q�}=kf�q�^a G�T,�h`ANtf�M�W�n?�Wh�������=�o<����E��a��3š�7u�>��Q�P{I1�1�ȍT����1``/P_����n�4R���ɚ8G��&NP#��a�߅�d���U}�Zy�o�۷��[�D8'
��`Y�������tC�t���=4t�>g�����<�f���-��@&�h�a�]�Թ��$�A�n�o��3ݡ|�M�9�RKѣ�}Sm�	uA^¯�f5k�J
d��9�yx�b\�.�0b�k�#��w�Nf���VУxjt�վd�C{  �_]��h=���S��b���ӌ�A�,�o��,�H�c��[(��s�TF&�����x������+P�* ����N\M�R;�S�V~<y�!�����F����X:}��^2����
�U�����H���O�:FwiuC���
����c����c�8ZX1Sk�`�Z��S-�v��	�-q�J��Ax:Q
dڃ�O�1P~p]s�2��{���9���q�@�0�� iM���o [ԁ8�{�I�o��΃l��'�i��������^���P	zbs5�Hx�q�� ������]��yk�h��T_q���Z���7Ja3��ѵV���\q������
�ͦ�?�:��'���6���IC)/�=�'�3$�����9.�dl�}��{DBZ�=�'��m�O1�I٪�q����I�i�XM����K�^�H�g�Ŋ�	��h���i�Ǭ��)�,ɀ#�	z�d!�x4	0���1n��A����ʙ�Åz�6�mq�`7�m	+T;@�ɾ�ǎ(�nɥ�'n-_�2j6��m�	��b�� ��V�|I���Z���_�C;�l�ޮ�7�~L8�F�2P�#ؘ;�A�^{��'����y��ٮMveU�ʨo�Z~禽�+&0N���L����˄3�z�t� �(��_�  ��[�^�-G�q^��uG�z����y�Vb���D������f4�x�6� A��r����0�=���+l4&je��DwJ��s�s�?�.��υ�7�� ���0��S|�%�����?�pJ `���8Цm�~�[.>��5YV��+��X����ڳz���"48�02�Oy~��l��L�p�A���=�2ƻm�4v�pi����r�PY������x�m��4w���_ +������ڨ�g �4*�)�����%��%��G
��$1'!�E�k���v��,�>��E��D�P���ܖ8#l�Ѽ�zҰ4��[���KYM+�#���&-̪O�#���Cc���GlV� "����!�i�>}��<"~`x�{v��=M�B�^�����
�D�ntH:����F"�)|��Rd�8Ub��O�:H:	�\�$��9Wr
�����Q�����M���U�5͂����L8*W����Q�M�<s+�h������\	pҟ�6>Z6P�#��q��t�i�@hkC�D��{�\&E�����o�],\��7�	1�k#��=�Xsf!܏tx�d@���_1��a7���	�{��=�Rx�~d��hu�� PE��eqc�����[68��/�S�GG�r���ް�*a��R��]�s�Y�8�1��
�/�H���)�B#u�e?0�S��
X%&��/�U�-F���'��g\a���C���#+?�gк����/IX�R�a�e��X�9i'��%�&��9��i�����j�ƹ��I	�+���+}X4vM/E"ur))T�>ꤡsuN�|!'�<��Kn�_�����F�mNʁ)��-�q���1�6��=�H��M;�t��U�����w����"	{�i�D�H�pՑ�k�ƽ�jk٢�d�]'R�k���D���gp�\t@z���XDGK au5�vYw�D��s�M������<�H��&���	0ˢ��av@V�I�����#�W>m�}����\��)i�8{�`[g��G��J�9}V۱��{�ܴ��ӚԬB��~��y�{}��f����B���D���&��A��_�B&Hx��vDK�r�H����{�G'0��=��H�����ReoK~�5��§9kҺ9��g@#S���G���2�:Viĳ�ύ
>l�H/�=�tM«�Fұ�ٛ����.�@���kmC�u��������M$���1���,ɾ��#�4њƊy�v2���b��m?5�y�}~�T�"Z�*P��
�s7��[p!f�=g�韲N�B�����	Cv�&輺Z	�Y�]Ļ+r�s�`������EZ�٣�'	|0;H�W��h#@�BnЭ��}T%�t�h�s��H0,y���wC��L|ͅN�=1p9�J�z�b��>BoX��b��Z��'��p�������
���Z1��4��{Y��f6u��H��q̃Sj���#Y�Y�x��*cA�J)tU�(׻+�nG�h�"��Ks"��-5�#"�7T1�u�AvZ���_���M-��ش�ό:.�~�,l������v�vqmߠ����F4��>�&��Y_x^��I"r]z#@Cr�N=L��Ս+����z�6���Mp4Bo1n��v��p�/�-IP�u,���m��wU�<\j���=ҋ�/��R�>�K���B��P���ܧ6�[��1[�������ϗ�G�{�*��yx����쮖Q�Q����6H�ʇ
�Ӻ�)��Ά`�8AP�<U�%G-˂�0���7H0�Yk�P��z��j�̈́��P�On[S�ݺ5�	�R:���
񅢽�������&��=��S<���.'*s�Ϸ�I���HdU��
:C@���Ғ��Uग�|�$�ٙ*$e��*��@#a��-����.u�'��gJ3��5V��r������H6�@BI�D���"�i�)h���N[�6xY���b	<�6ϗ^g��e|�t���	jQkm&H�7�η��y�MWm�&��>Pņ*����:�CY_?ߓ�UA��I�2��kh��&W}$!h���L�S7�\�Nk���Z 8��d�9����חr�ո����T�	��r���Y@?O�S�>9��#�oj�-�I�5-�Iؾi��wDf���6���U�}P%��_�yVn�����4�s�M:r]�#�K��`�$���Rg�m�en�E�@j�`a�{Y�n�Hq6��`�v%�!溴���\�Ǐh�|H�*�<�f�ApqV`ȇ�ё'Q�1����n�wB-Y������1�q�Og�]&�H�����
U3���s�6d�W�A�P�?B���m�55F������VY�)ޘ�V�LD��1���)+��=��G�Dcxg�?Q�	����ũfVp��W)���A%��-{O��\:����y������u�3��[��s�/���b����r�eZ��8�������E�0a�c�	P��-%N%G���!ԟ���[7bV��aC����=���$��c�C[d�>�[���%��|���Cd�Wn�Q�~�W�鋨�?m6��I�� ֫J�W�L �����B��l��n�[Y��D,}��F�-�I1���r�slm��u���߲�#�6�����,�c�$_�iE��2��A'eݚ���Ivgۺ�P��_.jc�ax��� �,�6�"̆=vv���J�>ˮ�Oi�)b8���T�o̙�V�Wy���7�-�&j�����?"%
�2fR����@{�C�L�3�]u�8�"O���~Zx�f13��XT�w6�~ÒG�̩�_�>,4�N"-4�um�1���C���7�cR~�ZiX<X.���Ւ}����Z�6���a ���b�i�5���0�ର}�����^D���`�r�0o��e�=����	i�,!YT~Gح3'�ऒ;�W�fCj�T�Ww�0��6mz�`�����z��s$��vWJ�Sɖ�^t��Ĭ2�yba>й���/�h���?|b���¶7��6�[H.ʌ��٢uӝ
��vQ���g{���_���l"�^$�p}Gq�\�j�Ҍ0H&�Gr��\�a�8A���XҠe�:Y�3O�?�7N���Lц���%�`S�6=m^� loJ�оQ�@CZB�j��K����cN�^����hN������k5�x����yH.~�0#��>6^�����߉p�})*_
�g����ܒ����u|G�����$L����;�aR�E_����G[H��P�WL!�]�8�j��x ���H��O �.g4F�#"�-�t��,b�tM0�Nè�c��f;�i�5��l�Eg�a��Ȟ�h���`Uӽ���7�Le��b�OE#�GJ��ʌ���fǌ�,�ن������k��ߥ�%��ͱE�;�`�y���S�]���qmA�4�B��2�Y��MK�R���p� nq�4��($����XT04���	PS
�C0`ǯ��$_�gU`��9˼0���v.��O�IĽpy�d$��?� @�q����j޻�As-W�ub�ț�{�%!s�*���^6�E\N�"�>��'��	v���{��oX����bn��M��<�>j�/?X��������l�LW^��8�?/�Y�zZ�P���፨-a��b>z54���� �	�sXd��������e�D�"��!�!+/�Ϟ�AU�&k���"xGx&=�K7I�=�d��ĵoz���܍ /�����v(�Ν�2�b�3za�Y��
IW��2bbE!�.X�gH���v/���̯��#��y�ˈ,d����6��$��%Ԧ����! �N���t �Yx�l*�F�E��a��1��c?�E���I��%c���o$������ett]�~Jg�ho+`�e\F�]����b�u���,�k�١i�Z�0U��"ܱ�V]�������R��B|�~����T�G_w�4F�)�G�����ṑM�VJ5�2�IIvjNx��y88	D�S�7�~��0�H{��_!i�ܕ��{���2ph��z�-1`�<F��Irq�]	o͏$/�Y�	{�C�5�N�;ʌ@İ����,���I��Jj{�f�jPJ��v�]���1�k�@F�!��AU<��N*`+�!�����Z�#��m/q����#G��WO��"��Do7������3�R�#G�^�*�	���SkeSQֿ�a��%=y��p����*�#��|%�*~��ͤ6,�(�+d���2�;�����\�X��S�q�P�<����7̻�F��r�t���#U(��<��^�����p�E���C�A]�z���$:�RI�uRp@{MA.l+}d�١�P�KՄ�Po��!4ZI���	�Z&�\[�ѝ^

u����5��M���ߟM6-L�.*,����~��`3G(�1H���="�)�֫��̛�X�r{04:=맕�E_إ�x)ȭ�~cu�
���s��7<��M��zfp(�oL��7c�ú�D"likK�?x7,ޝfV?ȶ�;C��� ���&�;z[�gÿy������S�n�� 1 ��hꉱ�F)MZ��.�u1�I�9��w�p�] ]���6�i`v�3�rE��sV��O��`�)��Ǒ.l�	�,���+Cj$j����܉�����������$�;9jV縡�7�S��
O����>@�(�,lGu'���r$g��T81�V"��<�1}Y���{Ш�,u�����4��U�@���y��^`Hyɗǎj� -]J���p��
�w����l��#U�=��Y.E�gf������&
9�91pzCf��{J]܁���x�m�����
��2W����-�'��P�I{�����r�<J��0����ԵaB�X��	���5��
��\rĆ�m5Jw�WG�،hO��eG���F�q(4[҉��t(��9$璡��Τ��������=ר�r͟� ����Hȵ^��}=�1�h�py~�J��[��s���?����ja�H1oW���z~X�X�T��=�.0n*z��d����`o#oN��M�����ג60�ە����UE*�Q�2�^Pi�����(���O�O$�&�/Â�:0�F�J'����Kȇ�u+��x�Ԓ���@Y������ত�*ζ�eS����P��{Ǳ�"����^�mEt�D��� Z�X�ޯ-��.�S]�%�Ԩ�-t�w����W��W\�(�p�üv���_U���j�>���q͞+e)�\;y�.��m뚄��K��9�a�57�"D����G���Y�S�Z�r2dC��;x<��U8������Ӕ�������B��`YP�aP���7������`k~a��i��5��G١�������Q胇����M��.Y4Ĉ[������ܒnI$,g�1n����YP�ꝰ�oUU��}�LHMw"�	���\-E�Q�b������z� Ү	*�V�rB����A����t,ǉ��]�`+ʋ�GD��}�őrDI^��_u�_ ���C9���!5Ԍ'��,_|;Zl��Z�{�`�����R�韕mJ����yH�[x�kk�b�C��b6Y�֑��];n`�D@�&�j١L��t�����������$�;P�7�=Y�
5o+�Y\��� �}�v�#�9)ۃy�2��_4�/�6L�[��UJ�Y^�L��v�E�3�ᘷ����"�!~����LG&�1<����wh�>�6����6Au�Kqh3d��\xj���Ϲǒ�:
|kBX�I�E�vF��bF ח:y̩M�rw�V^j�� ��� �g�yO�����r/'����l[��i|�ǘn��~G��~���x��u:!9n��v �+��3T��3&��$�c�#�zhֆ�ECuG��ѡɢ�X�=q�u�}`�A�G EƁ�5Q}��JE�bc|��~�NS9�yjp��r�r������^���~����!'_�V�����U]fX��OF�g��J�[}�V����ټ��m%���X�z�tm��T4!��Ǖ�4w�6��*2��v�7�#�ʜYNA�t��Y���n�0e����3ѡ�~7�׹��!��gP��R�}0�fE�[�v�Z�\y�q1A�.28K,�����0.HqO��׬Ȍ�>�p��;�F�3#-�c��t,�x�(鶞�ȣ��s��)�%j�Ɓ�~�t��&���XK<(�5�/b��t�ц��'˞?�$rK�z�������g0�[+zn�ec���w���a���4�;&�G�T��ȷ~�o2�Ǥ�s&�w�0�y��݋�$�f�g�(&���t�������z�|�0��@���F���I��U��gt�+k��u9)o�g�du�mx�d�.)ɞ`���Ff]�Y��N��4/�ѯn����e1�J��FI%�_'��A��%av�]z{�2�o�_|N�Yt	C:�,��Ҕ`����<����dM n���`����L��R[@)k�3�M�����/Em�Ţ�j��lԋ��<�g3$�!e�:��\w]�K��5�$7�a��ClWk(L��ʰ�|i.'5C4��7a���o���;����K���-�e��3ÐWU3�8����v�|�\�æ�m4C����&���,�yDn�uk�Mu�,o�����y����N�MZQ,�œ�fD�q�`�^���W��8#�W��X��@��v��R�������^9X���d���vXZ\�N��H1���6��4�Ҳ�Z�6E�&Zbag�&���+�}f��m����C�y����=������7Gz�D�.�.���)܂�A�"��ꌟА�}�T:-�p��ů�v���.�[�Ot�q��@��\IH�@�5�(���CgA��2�o��
W�m9+.w��@�i���@@����j�ҟY�~�{��-��pE)��4����(c���3-"��I��X<]��_��J�a��*+��b��
�h�<���a�N��@lcx�Ҍo�*6����s0�t��H�9[�]��ʗ�gL��V6�N#�0����ŃA��~8��wֳ�tv���_Z����*	 ">J�e/|�nFoa ����#	N9/iv�x�V����D*|��s&��LL�3�]f�� ԯ�Z�,��'G�$�[,�c0���H\ij�/]"(��T: G�z�
�  ��T���
w���5����&:b�yE�0DC���nR̔R>�?�^Z�ӂ��'��-��F/�'8����IIQ��P;�3U��-m�wNg2q4�@kҎ.�U#�\�N,B?"���V�>�aj����-:j��0�����h�'P�yx	1�N�򮊖���pqX�&>�2n��Ό˔9rR�p��6)�[�s������~�y2��W��k�[	=�O�F W�}65ZѺ�����8 ��`y��Tt��2�l�`fPn���ت��ѿo<���Ŋ�ê���$�1��&��3�A�;�4~��i��m��!��dN�]1�lׇ����!�m�qU�5t�)�D.�N_֨���Bvhz�y�%9���!Z���ip�r�x��=L]
����Nnv���!OY�_�w�H-t���Q$�MQ���[cG(s�Co�=o��
g`Ntu��ɏ	^�L>������1��K���;����w�P^�}hS�ɑ��yZBv%���L�0+�|���ӼN���X��ț�st4y��/���MTؘ�ao�l�+���7."��b,1��S��4_�.���n-��{�5� r?3�3���>N�Z{��a=�)�R�]�E%V&�bn���!�VH���*����*ٹ��N˕2�t��
�
��m��SP��iY$R��<:4[���n���*�]���Z�x�WPl��5o9Νەi\M���M�c�����D���FF�v3�^��ܡ֨��
�C��]Qar�����
F���(M����9ۋб�D�x*�4H��;�]����I���|O�����ƿ�&���q���)�XD��mВ[yB7���j���V�@���2_o)����p����:��>�owK~��E���Tm�Be"AZ����,�峟i�kA��;s���IWc	�b��X��Uy
S�ޤ#�a����@���a �l1d�4���;T��ʪ��䐣��Ԓ$��@��t�̵,�<�ؒ�4Z� ��%��O��)�zG��N�vw�~�/8�응�8���@���l'�|Q"<25n���-�]u��ϋQJ��F�*�#�V'��Bt�{�RC8�]S�N�H��VG:��"~ȑ���|c_oJ�o�����o�l�me�r"����F�(7ݹ�r�Fݸ��c�)=+�7�b��1�_g�D�؂�Z�(
�֠�J
�
y��`���:�aAnZh~x,��&� ��)A�eW0�@.�o��	��aO���&.$*O�Dӟi�X�w̓�ұ��sa����K�0(�t��#�5�8#P����]����|�m�q}��:�)�d��?�ɪ����_ט��8���X�⵹�b�v|-{�
��w׮�ޒJ9h�;��j�*���n�,���ST����<SyZY��ƣ���$����P,�i�b|���)K����+D����6^ǭ�P�i�;)
O���:l��f��؜�3�|C��O]�,�6�$��$a�P�t���W�[����n���,�`&��7��Z�����ʖ]��*�i�|0(��>O��d�p.0l5�^�h�g�FB����#`�w�8Mc���Y޽,��8k����4����[�#;�����������~��9Rƭ�$��U?��ﱵO7bp>�~
���i��w"��ژ���`����rv��RI�q��Pm�Qr� �i(��v���W%#�1/UY��ҹa+'O�����E��k�U�"j����ˢ��dy�&�YY�p?4��[>�O��XG
KT�s]�W'N����x(b{���׏��t+��-$s(����%'�!�c����s��3���h8����C<�f]����u؅r��s���z�&�	�l�I�s�� ����س���.����c�eY�V��.�*Z��z�ҟ�ˉu���3��{w���pj]��+9�c�[({o�?��/�B����]m<ʷ��؟�����ҭ��xX����r-�׸ �F���T�ɗ����~�y$����ܶ�a͐+��`��
��ãb-v�!=�:�-�C8�Xu��j��	2մ �_�#��sY�ׇA��2O
�qKz�(�5���<�B4�[\_D�W$s�0�@�)����4=�A����~j%c��R8�奺��3���]�w�`=ao-Yn�=��ؾ���.S{�?���H+����ȝl����\��/Y��5�o������P��S<F`rz��Hvv�p!�dj�y�V4�W�X��[�Z�������~��q�|/w��Z��s�3��J0_�h�q��h\k�i�j���wh����Ǟ�E˴sn��T�Z��(�C�x��#!��+H�/Y6f�s�PG��E�J,ٵ�%Y{���'�,��	��EB�rٛ��o��Cv�R:-�)��Ve�!;�~ជP�(��o"�Y?�E��o)q����� ��hks�L��0�'�a�܃�YG#X�+]{��U���nNW�$�jxŶ�VTjgFm�����W!K�t��8�}]k�舵!A5�Ԣ7�A?F]�J/=��c"���@������a,q�8��a�`uO0�
�iԲ&�\p����6�Z/ǄksF�oe`��*�׹�I��d��]7��kK�3��ga�qV;���>v虚��ܢ���^Xǌt�0����t����a���#���;��r��>�!��; ��9�2��ե���U�i�N�hF�a"� �T���qac3@��u���j���_6���%�̺�����
�����1���D�U�Hܻ.��B��B�Ĉ��������ko䠥$�$�B����i���H��+�GW/����ډn�SI�B�O���������Qj�2ӔV��m���n����|\������sJd���Ʒ�Z����4�����u�;��֨�����sN��8B�(HKRmuZ<����"��=4������}�U$�1Q\�Cc�b�	$@o�Jo�ף��c��/ܧ�ӹ(&g�䋷ң����˹�
P�e�6⃟� �?hZoq��2[o�F�9łqr��!�&���sq�ҕu� p��c�;�\0��aA��<�V��ʀKy]ͱ��z��t5˩WdkO��������@p�6uX� ��ɸ �Oe �� J��Rjw.����F�%��3�C<z���y�-CwY�
��zM�pr�=r�{�]�aQ�� �i�Z���{M�ш�����_����2r��܏²�tr�18�r(���8f�l����r�j 4=S���ܮ�����U����
�����%
��v��C?�.�F$��`Kr��-&O�P
`��cTӠ�,;a\�ꗭ���\��ʩ�Ց�g?��v�#>x������Eq�����d�qR���;�8�߼&�v�]�k��Vb��G-<��)�c?�{E����ӯ#�"tg!����~R����h�2m��R�����ޯc��4{h�=xn.�N\5�4�����e�ۈp�'��FZF�͝X!��L����ޝ�C�Lx�W�@����P|��g ���@�: �)_�nA2����Mnj7j�R�
��+�F�{Ԛ�$�%��>$H����3�)($���u����n�43e�I�h���2-�R�t%] �n94��C(Y�H�C���[�sJ����Vh ؛*$��Yr`�	KgXFX��Nx����Όx�0k���Ba�����{s��\\�<
���!2���k̈́oЀ;���Eނ��N*�)�t��R��iv�'����qѵ�#��AK�ml	Ay*�A��m]ؒ6i����I~�7�p����8��{�% ;y"�wC��dM�����vl�f�j��o0f,|�!��:E ]����ɾ�F����}�B�.�'�A�!��RO�HD"����~��%g�Oa�J�˓�2��;{��m�_��P&�b�bff�]o�6�֦�L;We����x!-,>��F����K\+I��9WY�բ�)�{�Bey��	�f�9v&	�j9s)��[A7-Q��. �`�b��ϳ�4���2�*�a㰎QX��ꎵ�ц�����hA^sQN^�*�قOMZ����hw/��Z��qM[Q�)�=H����
���2z�y.�+��A�}?!,�v�Q��i��H���-���Sq��!/dӡ�v�������*���}$�*�3�3��_���@�ė�m�Y��d�P*�BhL@kBz��N~�P���?)O��cU���EM����8a�bI�6���W�݆+-���$���^Kd��]�T�m�I%&�~��/Ϻ�ʘ[�YZ�|��.��H7�t�G�;�"1���r���=��c��9j]`��<���x �n�ϝ꠪�c�{�>�O�����$Z�zD�������Ŵa�0��QcGd�gf �غ$Qb~Ξ@q�����
.��yh]!�s{���
C����A6�4�$��/���}����V�L^��߼���jE��Y���5�X{�6�k�n@��V?��۞��2:H߃�j<�8���!E-�&NJ� �z�}���QæE@��x7�!�B���-%�{�Cs��U��������#tj�젞��j��>3�Z^�d\	�F��v���k��"��YR`sD׏Ӛ����ɽ��|̡���(f�Ԑo�N���i��{�q�P��hQ���t��Ωv3�Dd��W/?��6�� �"&���88��ìk��:�Ҟ$�屢�$9i�[=(���t"�.3�ݑ��7k�@�Ol]j�^(]��{S��UV���=�7݃Mc��I�+f�vQlk_)�z}�6zHIkS���;dd}%�O���>��M
�D�m�����-)a2є����3� �`��N,��n��d����}N~u��ۛ��#��څ$���$j�		�A��{pd�GV��;�Ohz�/,#q����|�j��j��f�D����1���f�*+��i���ex�)�u�Nye���@�"�4��P6�����/�q�VF��
jF ׅWr�Dk��m-^��rx�4�0���ۮ�*	�N�^19�ɶ��h��vw�r�е�����5AM�e����Ų$)�������+���$�m���˺��*���S���z�a��Z_�.��v���d�����$�ʇ����S�ƽ� ̚ٛw�<�Yծ�a;gF�`&�1�
�ە&�vQl��f�6�?M;�5ٖdϒԜ-�l�j'n�Uŗ�-5%D��(,32�.�
�zUa��t���M��i\,���^ȝ���t�\P�@�3_��m�9b�6ǵ���`�[`���x���p���g�#E���^�󤟛u����<:��9�ټ
`�O��tOx{�i� q�{��S9�n�Wr7��c[�qj�l�y �����������[6�Hi��kvl,��a�)˖[���y�V)��Cw+*q�W�Tz^��+h��-Y������= �JSǸU�}�:%!\/,�0�)�2���BĠ���+-&X��ul+�v�g�Qګ:@t��ߺčV���|
(bM^%#�K�ή�ZM[�u�n�e�%ƥ�C�|�۳[�sEdm�O\�ٜ���x:snIc�A3�Vx����j�J �ZC.y��`��-�쓗CX9���8}�2�|�I
�*�7)����A:��{�ZZ�V������f$ =�D����z�"��]����T�M�Ggςc͘�,�rc�E"a�S��Tr*�a�NՖҥ��e�"+�Pa���xF���
(1��?��C�C���>�|�Y��R��jK�GM~{�x�5��H��EKȇvA7m�l�	�b᧋��rrGy����f;�^�uwډ5J��.8+P5�� �^D�@C	�k��>!����>E���l��j(��PGSC0�!+�<�I���	�ٖMo��%�@2m�о�$�Yh��P��<��ed�:DǏȻTc�G��QP8w�����̲ܵg�[x�Ӑ�v�`�׏���Pڴ���G�6~b�TVz'��%��Ød�:=��"$�ŝ ?6~�H��q`�Bt���m�����ֱB2��XS�aJƞ�}I�URy$>-�������"mr�>ˤ�i�J!��ޛ��1�Y`�K~!�%1Xv�H�ڑN�K�u<�,(�S�ͪWw$
��JM�
���^���˫T�?{��O)D|	m����pi̎lF�H�s�[�u�%<hs����u�du�`�%.*r��z�~	3}>[Xթi~$��M��U�XkZX�r�ݴW
��M>������ӷ��i(���J.y�̳4�?+d�T�1Ȱ�usLŋO��`D�y��]h��N�U>�j{� �e��]a�b:P�l�P��+eTU%e�eq;��F�K��R��C�7bȭsR$I�����Dw��4�:�%C�K;�E��t��	�j{��у����4���E�Ly)`�1���i6P����~,%hu�C����P�jS��Ij��?��X��c�U@ǁ-C� �D�(���ɚ��X�%�U8���SD4��2�
����'Z(ƅ�0�p�Z��ڦB抌���b'��f�0~���˄s5���e�R��Ay����w�튝N��[��)�v��UV��V�!�~���3������
7\kj�[�H�]6$V�6�����Tݾ���\Ɏг
�:���FҪ?����0�s0��cC�b��(�>� 
�nQ�7ˉ �s[��4|�|�e0��J��~�娗w���"S�5��+�gR��e��f��SK� &��i������n�N������ԅ���$�����O��G�+���9���3z�bf8,�H����a�	�yo�d}^�;/5De�����3��r�<�����\�j"S7X�Ϩʛ�o�+�r�mjp�3�|�3�S68b�[���Tq�|�y�;t������f��tC]�Ldy�O��$8�r�� �mu�V˵	I��{eT;
��q�� �q�C��.p1'v�M��ϙvjS���2��&�n�%;Ğ�#RӻEds泿ԴP�MvH�iF���A��O�$hV��+�r@x(w;��Zػl�j���6ņ�ͱL�����ۿ��8�b�E1m�%S��=��=��iN�����q�"�����6�e���bI�Ş]�����d:��/������K�������ͷ+�ǽr�n��hd�ؔ�����:��8�\B�$iB0M%�䠒@=N��!6Y"/de��֯4�EU�6IC+#q+�b�o��\m���c����$�y:�H�dᣊS�/Q�� 
(�q[��j�O2jh��E�����)M�7�$g���%'�<�,G �fĢ'�Ձե��B�BW5����C�;���!I0��g�ћ��G����	@,�G8a�~;���"]�x죙@�,R�pt-�P�S��KN��ij>�>?c�9	�lvK\�[�X��J���1��VΔ �d�O�JhMbs�4��7�n�љ���0��p`(��.pgMR��Y݈�8�n4K���J���1A(`�a�r�e�(jo݁��q�x58�%��i�|���ug��A���(tT���ҥ�����#�#�.6���mM�u�Cֻ	��D�"� ?ނ��Ɔ��`��ޖ_A ��Z�Ehx͉�����q:�.��a�����i�-�é���R�]�D
f�����5-�Ķo�%p�O�Cf\�H��,�9B�¥o��.��_U�jwU!7�V������i����V��v^����l�!���ρ4(@�<�c>�0�ʻ��$���#$�TkܽI/,:=�2_�Saҋ����ҋ��J�gV��ـ�آ�v�m��P��3�-1�~�.��4=� (K���@9$�ڸ���D�����9<1�Q/��H'�B�X�+9tX?����%.���K`|/$7}$R�i����@dp5��Ehc��UW�ד;�E� ����z�]���9E!�hn�=��#67E�����(�;׌t���+U勉l���I[�v��a>��	�n��V=���5�~g�L���%�?Mõ2�-��]�y�VI����Q7 Z�&���N��
��E|!��F y��t9O� u���?�?��b��N��RdNt3�`�k�'2���B���1�o�[l���٫��W�o��@f69b�G�R�-����(P���3�b�Eٯ������6�-�~��a�6$:�G6�䀚oL��u#n��)��B�6�Jl����y���S5�d�����G��n���_�&�[���<9�A�g�a�ҕd�p!�q�I��o$�$S�JB�X�έ<c ��}��k_�;Fc�ٚ�F��Ĝ�ʫf�x�����sJ��w�B�}9huu �*:� �?���1j����]a�Ud�1�/���������4t�d,��%,��c]��=.j
-����]�R2%��T��_�#�[\^����̼jvR��~���{~�?���'Y��0�bq}Xxl�^ע{5K�1_ս�-vc|�[��,���g�Dş~��M����7�a=rp9��<OY(�oxa����Ǎ�:3s����C؍��Au=k�ל/c*$H��8����[���1|{�:iYx��\B,�k�.l�RD�nIlWu-#-
�vjI�����"fr������1��Ɣ�f�߳�%��G��)U�����1s�i�kwu��\��[���Wf��5=-�U1q��y��M�h����hQ�,����E�=��/ ^���^���Ojd%5�V�`�M��M��H�x)��O��CrN64�����dő�Ō��R�F(E��u�S�i�l"�_����F��0�gQ���\1}m���
w�<'V��ǆ�>)�g1���y���}O���`#]a�G!E[Ja�{�i�D�	�	�pv�J��o����R�Ѷ��{�EV@[ǠA�;;c(���,p�V�$6���C6���o*(��"r-!G�����x�N�D1V[u��
�՚�jϋ�,*!��,P�>���s���4U� �o�vu���s!�]>��H
n��ʱ��%uV`0��t�Z'gQ�w/������SJ����+��kb½v����5�!<�+$L���Z��~w-'l�N�/�^p��"�N>}���·�H���&0nܼ��T s0v�NԎ���;��̕�X��BŹ�k��#M�o�mg�x^m�0S���8M����K���_�L ��N�ABTr#�e�R�B���>���щ���):�-ox����:��Q��=�l�C<9ʌ_������2&F����0�ƫ J*��C&&�z��=榚\(�g����s�
�Y���`Q�7U�ĞhC��b�̯��,�߼D#����1����<Ճ`�.zI�:�}5���9�f�v���-Y��䀽MJ��Y�)up,�$��RVI���ߍ5	��|9��Q"��[_�����l�4T�s��<f��Oib�V�" κ�h�6^���z��ޥ�����g��t�҂c���ޭ{��#�Ql��lo��c����q���g�
 ���_�X�T�P��=�HnO[S���|F�)�V��(�"K��N��\�|S�Z5}�+����xA�5{��E�C��\n��n�y�a?�	�OK3g��a�P�@�(6��Og� ��{v��UL���*�����;�ӱ��;�����Ӕ[@}z��I x�dS�e�'���ҝ�w�t��T��O��q~-~m��r�c���f�٢����P�����2�\e^�4��9m�AL�\(m�nR=|�گ F�܀-�j/��)[3��������Tk�O�g�r�+^�Mٚ�cJ��3�P+���T��<#j������+�5nĘ���S���Ê�.S7��b����Q
���S��:;V=���l�U|����,M�u����m۪�d�Dh�3�b;�;�^#Iho�y���Q���^�8�A�ՙ��:ܺ~���=�L����x�d�������]� kK�(��]�BG�ލΎ�u���ZF���t�����]'��S�w�Z܀���T[���wv=�j�	kU��T�5R(�%:T6�[�g��i���J�����R�=V"B<�}Χ�.�:!�Ȉ���	*ٶ�)jt�"u�H���K�w½��-N9r�vI)^B�s�V�Tyc?�	v�hc�������<�;���K�B�U�������cs����b ��P��cp��=��<|>`O��+Y��&������5����'�H�Vn��p^ZT���L�����0U
�=�D�2,-US���{�?�z��Cs�0�@s$/Է�R|�}TP�F�9�t��^��Ys���yQʠ�����+�3"�A�2!D���bUd�w���R���㣝�5��{��r������f����7�s�Qݏ���c�Y��.����/֡(N�O�����I/���y�ߛV&v|Z3x��N���������(p��M��A`(j"�P5�U��Q
I�a����r���LX+���z�؏x&�B��B[�<��^v�d�r3�_n����.�t��wu]��^�x!�dZ��W3$�Y#�u��/$�z�
E�{+8���'d��������+Q
wCj��D���.�Sg�P9�8&q����f�x� ;<��_����
�+�6��D���9��C����X�W� wGӤ��z�	��*Q�*�zJ}Jzxq��_U�5TKx����Oveꌇ�m?�|sJoUd��j�1T Џ���c�Q��-T��Ć=P$$�򼏨onz۲Z�s�.^�W��Ïa�o�C�Ҷq�EK̚��Q�"����7�����'c�F����.-]T�RN)�!e�7Y���P���-�k�����,s-L`+^~�x�O��%3���:��vrl[/M����rY��b���8e��?���9�����(�:HdF'7����6�P"3���n�1f��}���@���6�/9Ȗ��\t:.о�g�F��-Sd�&1A�)ѿ]��4>�K��㍜Ρ(մ�������M��=�VP3�U�a�(���*���EB�v��:����p�KT�i��\�7�ކ�V��M1�>A62�| :U�L0o�\���B�e7'g���d���[�o(܎�I=�q��� �^~\��?�����~$X�0�r�}2�c�[�79��8���<(@�k���p�}m�:��#g�H��I�]�Nde���~���*�{�?��4^�PD"1\��QY�޷���j>�X��m�{�u���rkE��^}c�D�jU��z����5vGɣ�7_��1U�fn��ҥ�#���ye>�~{
d�/� �LX5�6�Q*��c��h�ph��� �E`0���p|:Y��K��D��AUw*�6ƿ�R�ԥK�˪��Û�N���j'�e8t��Zb`�,�͠+����tN�R��/�u3�R�葍v�@�y(�Tm��	���a!�]@�V���Ǩ7x�9�r���Ꮊ|5���]J%��]j��Y�7P���'s�n�Cs;Qva��Z�0�
��D^�f�t1�T0�W�OtQ$g�Z��^t�[�*����3Ug3}�n�(4m�$s�[j����3��I'ZU��gUm����@��1���e�"$y�ƈZ�r@Z*�A���^(&ݩ|��ЁN�,Y��f�&�iΪ� LD9�c�g��e5'������]97�|�n�BM&��ec�a#��ߟ�rJ��u�䀽�zem�$W񉺁N���e���������Ųy|B�P��o�DD�#��w������I��c�5t��)���C�m��]0��Q��H�� Hk$�͗B��g�͢���}��Q�������M�����0bݐ�p�ҳ$oI&�]���ڕd` 䪰ù�	����*D�?�c-�j�ςO��}�P���ԧP�0��QDRi������E��Hrkj�[r��s�֯5c��u�r�^��;�<��@�B��x��٩�`f�)�yM�#���N#���y>���Z��=���l0�A�mU� ��Cvn��B!gJ\\kwV�n��y�� )|r�=��(�lw=d�u?/�p*�51(�җַq�����~OY�5����"�RX'�AAd�`��(�d��o�1�6�BA�K��U�]i�3j-黜�ӬIR�����#��ˑ�������2��P[�y����_-�в�B3�n��r�H�	�M�W �g*on����.c�J���1��N���p�����D{{/jq��AH5��/Y�,�1��ӓ�&mMd�.��8X���l��(��'q.�f(���] ?��9���Ur�;(�
"�l�eq�,��������6�U�8�:vR\&�?l �H���_���8P7���Ib�KEF�w�����W1椢�a}n�?j�w�&����EՈj�SSP3�yT҆����7	遏� w`�(;�-�G&ZG��� i��ӌ�֮��;���2�ٗ瞃�"%i��\��<�{���]�2g��E�O8��v�|�,}�t?�U����D<�@���`g�[�n���	y)�d����6/]���������Ul�Sc�Z�1����c��=��<��P*r��ޖc�x�o�׍��SO�OZ�60y��ns�)Z�	�l·*^�w�j���MC�d�� ����Iz�<$�7����	��+�$�]:����q��_�s.j��M@�	���7�k�C#�xC��3���c$�>z���T�!C��t������
 ��Ɂx,��	�oٮe��}���{�>�n@Kk���nW�F?�O���0GEۈ��������M���h�-0�fI��K4Ι�@�
EIT��{���l�fԅӺBeT�:������{�l�X����$~����b�� �g�\�^�Xz7�>��[_��B�Q.�UC%�YK(��T=�������^�L��B�W$F��|��}����3ҥĿ��_�j���ȱaH❓F��!�-Fu��"<j-���r}4�[�wT XnQV;�i6�XaR�n��EG$a� m��UM��][�(���X�Q/�6*,U�/a�;r�'�8vī��SyTг�V$L���w1�3���D�����n��7ص(g�����^��j�����^dQHEw+�3�x�.t�q��bM�n�6�=a:G���D݌ۖ�%U>�ոn��Vێz'F��\[���k�mhlb�2��j*I0\��F��+ΤUr���䌬�-u�pU�L}Ët�g{��IZ��T�<(�[��.�|+����Ώ_f���)d�l���1��~ɫ��i���aBlS,હ)I�W/�Ō+8B�T|��}:��U��}TPx|�E[����[�1)�z>�Y�f��Ԉ����{B:V����
�
	奖f��w5�f��rIP�;���#o6e�:v�{�P�P���FI�	K(�\�W15�b�Z���ʎi�b��s��I���X�s�����{<�>���Y�mh[��K9`���B�*�z��n_�DQJ{O2��ku����]`H�5x��z��-q@Cn��:>#�D(Ɔ:�(e�E�)�Ѹ}F\S����n9�!}�����k�r�pД�5��;��2��"u`(��^��7�V��&��#!�$}�o�Ai�5|�!,�Ö�ʹf=��� Q���f����h5�����G�yA~����u�(�Si�֍=@E׳�+�7<��V¢�g\F�͛GpZ(/�f����(ߧ9�.ܡ��}���i�G�#�'��	��[���LTȦ�Z��{�lU"�{+a��S�)s|nƌ1����w7�����*�vY�L��iFDl��>k���������ڮ0�u׵���3~�{�l���ѯ�߬��NE��Szg#p(M��u:4���F�ܕ�"�T�6}`��7M�W�Ԗ����H�7f�z�v��C�B�g�/%S�J�1�n�-�w����к�Y��t��^	N���f��N�t�A	�W��6��S��5H8m�>�4U��d���h��94�!sۨ�TtD_/�a����$�OELRXO����~@$�.��9d���(� p&�2�:�w�}8T�Ĳ2��:��ށ97D���@�N����������$u&1�$~i�ˆiη>On�Fi�MM�w����q7;�6iy�R�?�w��K�-K��KeCc�������-_\��F��Q��|�Y��Fc���jK�M+iRV��f��C�}�"�V�{�p)Vs��ŭ�;,nf�(N 
���4��u8̄����]X���#�I�3�B�4��b�V�\E�����pz���2��,�+���[��\^�5�������Ժb	�m�I0d���K{�G�aL�S&�*2��2ث"<�B ���zdO�>o�y�=K�B�[�cjz���,�����e��7ڠe�����/�����W�6NTi�q%����_��ľQ@����zE(�f��H�d��%�Sj�v�y,	^V�m̢w�M��˛��.���4F�F_#�#%ў8R/E� �1g�LY�i[틿ڦy<@��7I�4��9�Y�Z%ᗵ������¼P��V��V(>� ��I�k���D:�� d��U�_	���)G�Rn��b�O<�Y/�E&fڙ�ݦp4�?��'�B�z�*${qX��|���.� �?�)gsj��IK���ō�.��@�h��G��N��at���a�3�^J���.���$������m*���!��8AUu!{���r�D�wa:Wx�p^b�}�H��;
`�i�BR(�K3��q*�AT�͛��	�V�����j�kBaq��P/�6���	�a+Â�Q�� s�����������-���B-F�[b��L����V���#$ ��A��ѻ�q��mA��ݢq���=�_�Z)�X��r�`�̥�ÀEG�}9RM��~���V�F�b��9��4�ab� ʬ�7��ҹ�6(�d�Mk
��M�?�5M��
�4�B-~�n&*��D�7HǊSpϊ�%e�L�:��dd� ~3�%UΜ�<u!_I��ĪkI�ָ����߄g��+�l�r��x'R���=�b�r�B�e�]��C
ì5�a�9�5PA�A b (�o���֡��N��%�/��[��>���R���u"qp8|���o��p9�C:/MJ2�(�(�Ud���0��Ql��"���9m��i��\~��#N�7����(�q6�?��lWb�a8�`mm~/�C���<��X��2�#�r����fS�J;U