--megafunction wizard: %Altera SOPC Builder%
--GENERATION: STANDARD
--VERSION: WM1.0


--Legal Notice: (C)2013 Altera Corporation. All rights reserved.  Your
--use of Altera Corporation's design tools, logic functions and other
--software and tools, and its AMPP partner logic functions, and any
--output files any of the foregoing (including device programming or
--simulation files), and any associated documentation or information are
--expressly subject to the terms and conditions of the Altera Program
--License Subscription Agreement or other applicable license agreement,
--including, without limitation, that your use is for the sole purpose
--of programming logic devices manufactured by Altera and sold by Altera
--or its authorized distributors.  Please refer to the applicable
--agreement for further details.


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity dipsw_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal dipsw_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                 signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                 signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read : IN STD_LOGIC;
                 signal peripheral_bridge_m1_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_dipsw_s1_end_xfer : OUT STD_LOGIC;
                 signal dipsw_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal dipsw_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal dipsw_s1_reset_n : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_granted_dipsw_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_dipsw_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_dipsw_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_requests_dipsw_s1 : OUT STD_LOGIC
              );
end entity dipsw_s1_arbitrator;


architecture europa of dipsw_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal dipsw_s1_allgrants :  STD_LOGIC;
                signal dipsw_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal dipsw_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal dipsw_s1_any_continuerequest :  STD_LOGIC;
                signal dipsw_s1_arb_counter_enable :  STD_LOGIC;
                signal dipsw_s1_arb_share_counter :  STD_LOGIC;
                signal dipsw_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal dipsw_s1_arb_share_set_values :  STD_LOGIC;
                signal dipsw_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal dipsw_s1_begins_xfer :  STD_LOGIC;
                signal dipsw_s1_end_xfer :  STD_LOGIC;
                signal dipsw_s1_firsttransfer :  STD_LOGIC;
                signal dipsw_s1_grant_vector :  STD_LOGIC;
                signal dipsw_s1_in_a_read_cycle :  STD_LOGIC;
                signal dipsw_s1_in_a_write_cycle :  STD_LOGIC;
                signal dipsw_s1_master_qreq_vector :  STD_LOGIC;
                signal dipsw_s1_non_bursting_master_requests :  STD_LOGIC;
                signal dipsw_s1_reg_firsttransfer :  STD_LOGIC;
                signal dipsw_s1_slavearbiterlockenable :  STD_LOGIC;
                signal dipsw_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal dipsw_s1_unreg_firsttransfer :  STD_LOGIC;
                signal dipsw_s1_waits_for_read :  STD_LOGIC;
                signal dipsw_s1_waits_for_write :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_dipsw_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_granted_dipsw_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_qualified_request_dipsw_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_requests_dipsw_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal peripheral_bridge_m1_continuerequest :  STD_LOGIC;
                signal peripheral_bridge_m1_saved_grant_dipsw_s1 :  STD_LOGIC;
                signal shifted_address_to_dipsw_s1_from_peripheral_bridge_m1 :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal wait_for_dipsw_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT dipsw_s1_end_xfer;
    end if;

  end process;

  dipsw_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_peripheral_bridge_m1_qualified_request_dipsw_s1);
  --assign dipsw_s1_readdata_from_sa = dipsw_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  dipsw_s1_readdata_from_sa <= dipsw_s1_readdata;
  internal_peripheral_bridge_m1_requests_dipsw_s1 <= ((to_std_logic(((Std_Logic_Vector'(peripheral_bridge_m1_address_to_slave(12 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("0001001100000")))) AND peripheral_bridge_m1_chipselect)) AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --dipsw_s1_arb_share_counter set values, which is an e_mux
  dipsw_s1_arb_share_set_values <= std_logic'('1');
  --dipsw_s1_non_bursting_master_requests mux, which is an e_mux
  dipsw_s1_non_bursting_master_requests <= internal_peripheral_bridge_m1_requests_dipsw_s1;
  --dipsw_s1_any_bursting_master_saved_grant mux, which is an e_mux
  dipsw_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --dipsw_s1_arb_share_counter_next_value assignment, which is an e_assign
  dipsw_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(dipsw_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(dipsw_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(dipsw_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(dipsw_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --dipsw_s1_allgrants all slave grants, which is an e_mux
  dipsw_s1_allgrants <= dipsw_s1_grant_vector;
  --dipsw_s1_end_xfer assignment, which is an e_assign
  dipsw_s1_end_xfer <= NOT ((dipsw_s1_waits_for_read OR dipsw_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_dipsw_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_dipsw_s1 <= dipsw_s1_end_xfer AND (((NOT dipsw_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --dipsw_s1_arb_share_counter arbitration counter enable, which is an e_assign
  dipsw_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_dipsw_s1 AND dipsw_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_dipsw_s1 AND NOT dipsw_s1_non_bursting_master_requests));
  --dipsw_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dipsw_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(dipsw_s1_arb_counter_enable) = '1' then 
        dipsw_s1_arb_share_counter <= dipsw_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --dipsw_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dipsw_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((dipsw_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_dipsw_s1)) OR ((end_xfer_arb_share_counter_term_dipsw_s1 AND NOT dipsw_s1_non_bursting_master_requests)))) = '1' then 
        dipsw_s1_slavearbiterlockenable <= dipsw_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --peripheral_bridge/m1 dipsw/s1 arbiterlock, which is an e_assign
  peripheral_bridge_m1_arbiterlock <= dipsw_s1_slavearbiterlockenable AND peripheral_bridge_m1_continuerequest;
  --dipsw_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  dipsw_s1_slavearbiterlockenable2 <= dipsw_s1_arb_share_counter_next_value;
  --peripheral_bridge/m1 dipsw/s1 arbiterlock2, which is an e_assign
  peripheral_bridge_m1_arbiterlock2 <= dipsw_s1_slavearbiterlockenable2 AND peripheral_bridge_m1_continuerequest;
  --dipsw_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  dipsw_s1_any_continuerequest <= std_logic'('1');
  --peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  peripheral_bridge_m1_continuerequest <= std_logic'('1');
  internal_peripheral_bridge_m1_qualified_request_dipsw_s1 <= internal_peripheral_bridge_m1_requests_dipsw_s1 AND NOT ((((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid peripheral_bridge_m1_read_data_valid_dipsw_s1, which is an e_mux
  peripheral_bridge_m1_read_data_valid_dipsw_s1 <= (internal_peripheral_bridge_m1_granted_dipsw_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect))) AND NOT dipsw_s1_waits_for_read;
  --master is always granted when requested
  internal_peripheral_bridge_m1_granted_dipsw_s1 <= internal_peripheral_bridge_m1_qualified_request_dipsw_s1;
  --peripheral_bridge/m1 saved-grant dipsw/s1, which is an e_assign
  peripheral_bridge_m1_saved_grant_dipsw_s1 <= internal_peripheral_bridge_m1_requests_dipsw_s1;
  --allow new arb cycle for dipsw/s1, which is an e_assign
  dipsw_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  dipsw_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  dipsw_s1_master_qreq_vector <= std_logic'('1');
  --dipsw_s1_reset_n assignment, which is an e_assign
  dipsw_s1_reset_n <= reset_n;
  --dipsw_s1_firsttransfer first transaction, which is an e_assign
  dipsw_s1_firsttransfer <= A_WE_StdLogic((std_logic'(dipsw_s1_begins_xfer) = '1'), dipsw_s1_unreg_firsttransfer, dipsw_s1_reg_firsttransfer);
  --dipsw_s1_unreg_firsttransfer first transaction, which is an e_assign
  dipsw_s1_unreg_firsttransfer <= NOT ((dipsw_s1_slavearbiterlockenable AND dipsw_s1_any_continuerequest));
  --dipsw_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dipsw_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(dipsw_s1_begins_xfer) = '1' then 
        dipsw_s1_reg_firsttransfer <= dipsw_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --dipsw_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  dipsw_s1_beginbursttransfer_internal <= dipsw_s1_begins_xfer;
  shifted_address_to_dipsw_s1_from_peripheral_bridge_m1 <= peripheral_bridge_m1_address_to_slave;
  --dipsw_s1_address mux, which is an e_mux
  dipsw_s1_address <= A_EXT (A_SRL(shifted_address_to_dipsw_s1_from_peripheral_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_dipsw_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_dipsw_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_dipsw_s1_end_xfer <= dipsw_s1_end_xfer;
    end if;

  end process;

  --dipsw_s1_waits_for_read in a cycle, which is an e_mux
  dipsw_s1_waits_for_read <= dipsw_s1_in_a_read_cycle AND dipsw_s1_begins_xfer;
  --dipsw_s1_in_a_read_cycle assignment, which is an e_assign
  dipsw_s1_in_a_read_cycle <= internal_peripheral_bridge_m1_granted_dipsw_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= dipsw_s1_in_a_read_cycle;
  --dipsw_s1_waits_for_write in a cycle, which is an e_mux
  dipsw_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(dipsw_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --dipsw_s1_in_a_write_cycle assignment, which is an e_assign
  dipsw_s1_in_a_write_cycle <= internal_peripheral_bridge_m1_granted_dipsw_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= dipsw_s1_in_a_write_cycle;
  wait_for_dipsw_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  peripheral_bridge_m1_granted_dipsw_s1 <= internal_peripheral_bridge_m1_granted_dipsw_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_qualified_request_dipsw_s1 <= internal_peripheral_bridge_m1_qualified_request_dipsw_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_requests_dipsw_s1 <= internal_peripheral_bridge_m1_requests_dipsw_s1;
--synthesis translate_off
    --dipsw/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --peripheral_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_peripheral_bridge_m1_requests_dipsw_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line, now);
          write(write_line, string'(": "));
          write(write_line, string'("peripheral_bridge/m1 drove 0 on its 'burstcount' port while accessing slave dipsw/s1"));
          write(output, write_line.all);
          deallocate (write_line);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity gpio0_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal gpio0_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                 signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                 signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read : IN STD_LOGIC;
                 signal peripheral_bridge_m1_write : IN STD_LOGIC;
                 signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_gpio0_s1_end_xfer : OUT STD_LOGIC;
                 signal gpio0_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal gpio0_s1_chipselect : OUT STD_LOGIC;
                 signal gpio0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal gpio0_s1_reset_n : OUT STD_LOGIC;
                 signal gpio0_s1_write_n : OUT STD_LOGIC;
                 signal gpio0_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal peripheral_bridge_m1_granted_gpio0_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_gpio0_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_gpio0_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_requests_gpio0_s1 : OUT STD_LOGIC
              );
end entity gpio0_s1_arbitrator;


architecture europa of gpio0_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_gpio0_s1 :  STD_LOGIC;
                signal gpio0_s1_allgrants :  STD_LOGIC;
                signal gpio0_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal gpio0_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal gpio0_s1_any_continuerequest :  STD_LOGIC;
                signal gpio0_s1_arb_counter_enable :  STD_LOGIC;
                signal gpio0_s1_arb_share_counter :  STD_LOGIC;
                signal gpio0_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal gpio0_s1_arb_share_set_values :  STD_LOGIC;
                signal gpio0_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal gpio0_s1_begins_xfer :  STD_LOGIC;
                signal gpio0_s1_end_xfer :  STD_LOGIC;
                signal gpio0_s1_firsttransfer :  STD_LOGIC;
                signal gpio0_s1_grant_vector :  STD_LOGIC;
                signal gpio0_s1_in_a_read_cycle :  STD_LOGIC;
                signal gpio0_s1_in_a_write_cycle :  STD_LOGIC;
                signal gpio0_s1_master_qreq_vector :  STD_LOGIC;
                signal gpio0_s1_non_bursting_master_requests :  STD_LOGIC;
                signal gpio0_s1_reg_firsttransfer :  STD_LOGIC;
                signal gpio0_s1_slavearbiterlockenable :  STD_LOGIC;
                signal gpio0_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal gpio0_s1_unreg_firsttransfer :  STD_LOGIC;
                signal gpio0_s1_waits_for_read :  STD_LOGIC;
                signal gpio0_s1_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_granted_gpio0_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_qualified_request_gpio0_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_requests_gpio0_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal peripheral_bridge_m1_continuerequest :  STD_LOGIC;
                signal peripheral_bridge_m1_saved_grant_gpio0_s1 :  STD_LOGIC;
                signal shifted_address_to_gpio0_s1_from_peripheral_bridge_m1 :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal wait_for_gpio0_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT gpio0_s1_end_xfer;
    end if;

  end process;

  gpio0_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_peripheral_bridge_m1_qualified_request_gpio0_s1);
  --assign gpio0_s1_readdata_from_sa = gpio0_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  gpio0_s1_readdata_from_sa <= gpio0_s1_readdata;
  internal_peripheral_bridge_m1_requests_gpio0_s1 <= to_std_logic(((Std_Logic_Vector'(peripheral_bridge_m1_address_to_slave(12 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("0001010000000")))) AND peripheral_bridge_m1_chipselect;
  --gpio0_s1_arb_share_counter set values, which is an e_mux
  gpio0_s1_arb_share_set_values <= std_logic'('1');
  --gpio0_s1_non_bursting_master_requests mux, which is an e_mux
  gpio0_s1_non_bursting_master_requests <= internal_peripheral_bridge_m1_requests_gpio0_s1;
  --gpio0_s1_any_bursting_master_saved_grant mux, which is an e_mux
  gpio0_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --gpio0_s1_arb_share_counter_next_value assignment, which is an e_assign
  gpio0_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(gpio0_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpio0_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(gpio0_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpio0_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --gpio0_s1_allgrants all slave grants, which is an e_mux
  gpio0_s1_allgrants <= gpio0_s1_grant_vector;
  --gpio0_s1_end_xfer assignment, which is an e_assign
  gpio0_s1_end_xfer <= NOT ((gpio0_s1_waits_for_read OR gpio0_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_gpio0_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_gpio0_s1 <= gpio0_s1_end_xfer AND (((NOT gpio0_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --gpio0_s1_arb_share_counter arbitration counter enable, which is an e_assign
  gpio0_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_gpio0_s1 AND gpio0_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_gpio0_s1 AND NOT gpio0_s1_non_bursting_master_requests));
  --gpio0_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpio0_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(gpio0_s1_arb_counter_enable) = '1' then 
        gpio0_s1_arb_share_counter <= gpio0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --gpio0_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpio0_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((gpio0_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_gpio0_s1)) OR ((end_xfer_arb_share_counter_term_gpio0_s1 AND NOT gpio0_s1_non_bursting_master_requests)))) = '1' then 
        gpio0_s1_slavearbiterlockenable <= gpio0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --peripheral_bridge/m1 gpio0/s1 arbiterlock, which is an e_assign
  peripheral_bridge_m1_arbiterlock <= gpio0_s1_slavearbiterlockenable AND peripheral_bridge_m1_continuerequest;
  --gpio0_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  gpio0_s1_slavearbiterlockenable2 <= gpio0_s1_arb_share_counter_next_value;
  --peripheral_bridge/m1 gpio0/s1 arbiterlock2, which is an e_assign
  peripheral_bridge_m1_arbiterlock2 <= gpio0_s1_slavearbiterlockenable2 AND peripheral_bridge_m1_continuerequest;
  --gpio0_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  gpio0_s1_any_continuerequest <= std_logic'('1');
  --peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  peripheral_bridge_m1_continuerequest <= std_logic'('1');
  internal_peripheral_bridge_m1_qualified_request_gpio0_s1 <= internal_peripheral_bridge_m1_requests_gpio0_s1 AND NOT ((((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid peripheral_bridge_m1_read_data_valid_gpio0_s1, which is an e_mux
  peripheral_bridge_m1_read_data_valid_gpio0_s1 <= (internal_peripheral_bridge_m1_granted_gpio0_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect))) AND NOT gpio0_s1_waits_for_read;
  --gpio0_s1_writedata mux, which is an e_mux
  gpio0_s1_writedata <= peripheral_bridge_m1_writedata;
  --master is always granted when requested
  internal_peripheral_bridge_m1_granted_gpio0_s1 <= internal_peripheral_bridge_m1_qualified_request_gpio0_s1;
  --peripheral_bridge/m1 saved-grant gpio0/s1, which is an e_assign
  peripheral_bridge_m1_saved_grant_gpio0_s1 <= internal_peripheral_bridge_m1_requests_gpio0_s1;
  --allow new arb cycle for gpio0/s1, which is an e_assign
  gpio0_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  gpio0_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  gpio0_s1_master_qreq_vector <= std_logic'('1');
  --gpio0_s1_reset_n assignment, which is an e_assign
  gpio0_s1_reset_n <= reset_n;
  gpio0_s1_chipselect <= internal_peripheral_bridge_m1_granted_gpio0_s1;
  --gpio0_s1_firsttransfer first transaction, which is an e_assign
  gpio0_s1_firsttransfer <= A_WE_StdLogic((std_logic'(gpio0_s1_begins_xfer) = '1'), gpio0_s1_unreg_firsttransfer, gpio0_s1_reg_firsttransfer);
  --gpio0_s1_unreg_firsttransfer first transaction, which is an e_assign
  gpio0_s1_unreg_firsttransfer <= NOT ((gpio0_s1_slavearbiterlockenable AND gpio0_s1_any_continuerequest));
  --gpio0_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpio0_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(gpio0_s1_begins_xfer) = '1' then 
        gpio0_s1_reg_firsttransfer <= gpio0_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --gpio0_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  gpio0_s1_beginbursttransfer_internal <= gpio0_s1_begins_xfer;
  --~gpio0_s1_write_n assignment, which is an e_mux
  gpio0_s1_write_n <= NOT ((internal_peripheral_bridge_m1_granted_gpio0_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect))));
  shifted_address_to_gpio0_s1_from_peripheral_bridge_m1 <= peripheral_bridge_m1_address_to_slave;
  --gpio0_s1_address mux, which is an e_mux
  gpio0_s1_address <= A_EXT (A_SRL(shifted_address_to_gpio0_s1_from_peripheral_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_gpio0_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_gpio0_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_gpio0_s1_end_xfer <= gpio0_s1_end_xfer;
    end if;

  end process;

  --gpio0_s1_waits_for_read in a cycle, which is an e_mux
  gpio0_s1_waits_for_read <= gpio0_s1_in_a_read_cycle AND gpio0_s1_begins_xfer;
  --gpio0_s1_in_a_read_cycle assignment, which is an e_assign
  gpio0_s1_in_a_read_cycle <= internal_peripheral_bridge_m1_granted_gpio0_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= gpio0_s1_in_a_read_cycle;
  --gpio0_s1_waits_for_write in a cycle, which is an e_mux
  gpio0_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpio0_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --gpio0_s1_in_a_write_cycle assignment, which is an e_assign
  gpio0_s1_in_a_write_cycle <= internal_peripheral_bridge_m1_granted_gpio0_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= gpio0_s1_in_a_write_cycle;
  wait_for_gpio0_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  peripheral_bridge_m1_granted_gpio0_s1 <= internal_peripheral_bridge_m1_granted_gpio0_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_qualified_request_gpio0_s1 <= internal_peripheral_bridge_m1_qualified_request_gpio0_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_requests_gpio0_s1 <= internal_peripheral_bridge_m1_requests_gpio0_s1;
--synthesis translate_off
    --gpio0/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --peripheral_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line1 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_peripheral_bridge_m1_requests_gpio0_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line1, now);
          write(write_line1, string'(": "));
          write(write_line1, string'("peripheral_bridge/m1 drove 0 on its 'burstcount' port while accessing slave gpio0/s1"));
          write(output, write_line1.all);
          deallocate (write_line1);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ipl_memory_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal ipl_memory_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_6_downstream_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_burst_6_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_6_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_6_downstream_latency_counter : IN STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_7_downstream_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_burst_7_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_7_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_7_downstream_latency_counter : IN STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_ipl_memory_s1_end_xfer : OUT STD_LOGIC;
                 signal ipl_memory_s1_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal ipl_memory_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal ipl_memory_s1_chipselect : OUT STD_LOGIC;
                 signal ipl_memory_s1_clken : OUT STD_LOGIC;
                 signal ipl_memory_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ipl_memory_s1_reset : OUT STD_LOGIC;
                 signal ipl_memory_s1_write : OUT STD_LOGIC;
                 signal ipl_memory_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_requests_ipl_memory_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_granted_ipl_memory_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_requests_ipl_memory_s1 : OUT STD_LOGIC
              );
end entity ipl_memory_s1_arbitrator;


architecture europa of ipl_memory_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_ipl_memory_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_6_downstream_requests_ipl_memory_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_7_downstream_granted_ipl_memory_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_7_downstream_requests_ipl_memory_s1 :  STD_LOGIC;
                signal ipl_memory_s1_allgrants :  STD_LOGIC;
                signal ipl_memory_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal ipl_memory_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal ipl_memory_s1_any_continuerequest :  STD_LOGIC;
                signal ipl_memory_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ipl_memory_s1_arb_counter_enable :  STD_LOGIC;
                signal ipl_memory_s1_arb_share_counter :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ipl_memory_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ipl_memory_s1_arb_share_set_values :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ipl_memory_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ipl_memory_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal ipl_memory_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal ipl_memory_s1_begins_xfer :  STD_LOGIC;
                signal ipl_memory_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ipl_memory_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ipl_memory_s1_end_xfer :  STD_LOGIC;
                signal ipl_memory_s1_firsttransfer :  STD_LOGIC;
                signal ipl_memory_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ipl_memory_s1_in_a_read_cycle :  STD_LOGIC;
                signal ipl_memory_s1_in_a_write_cycle :  STD_LOGIC;
                signal ipl_memory_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ipl_memory_s1_non_bursting_master_requests :  STD_LOGIC;
                signal ipl_memory_s1_reg_firsttransfer :  STD_LOGIC;
                signal ipl_memory_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ipl_memory_s1_slavearbiterlockenable :  STD_LOGIC;
                signal ipl_memory_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal ipl_memory_s1_unreg_firsttransfer :  STD_LOGIC;
                signal ipl_memory_s1_waits_for_read :  STD_LOGIC;
                signal ipl_memory_s1_waits_for_write :  STD_LOGIC;
                signal last_cycle_nios2_fpu_burst_6_downstream_granted_slave_ipl_memory_s1 :  STD_LOGIC;
                signal last_cycle_nios2_fpu_burst_7_downstream_granted_slave_ipl_memory_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_arbiterlock :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_arbiterlock2 :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1_shift_register :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1_shift_register_in :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_saved_grant_ipl_memory_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_arbiterlock :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_arbiterlock2 :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1_shift_register :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1_shift_register_in :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_saved_grant_ipl_memory_s1 :  STD_LOGIC;
                signal p1_nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1_shift_register :  STD_LOGIC;
                signal p1_nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1_shift_register :  STD_LOGIC;
                signal shifted_address_to_ipl_memory_s1_from_nios2_fpu_burst_6_downstream :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal shifted_address_to_ipl_memory_s1_from_nios2_fpu_burst_7_downstream :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal wait_for_ipl_memory_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT ipl_memory_s1_end_xfer;
    end if;

  end process;

  ipl_memory_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1 OR internal_nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1));
  --assign ipl_memory_s1_readdata_from_sa = ipl_memory_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  ipl_memory_s1_readdata_from_sa <= ipl_memory_s1_readdata;
  internal_nios2_fpu_burst_6_downstream_requests_ipl_memory_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_6_downstream_read OR nios2_fpu_burst_6_downstream_write)))))));
  --ipl_memory_s1_arb_share_counter set values, which is an e_mux
  ipl_memory_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_6_downstream_granted_ipl_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_6_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_7_downstream_granted_ipl_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_7_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_6_downstream_granted_ipl_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_6_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_7_downstream_granted_ipl_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_7_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001"))))), 4);
  --ipl_memory_s1_non_bursting_master_requests mux, which is an e_mux
  ipl_memory_s1_non_bursting_master_requests <= std_logic'('0');
  --ipl_memory_s1_any_bursting_master_saved_grant mux, which is an e_mux
  ipl_memory_s1_any_bursting_master_saved_grant <= ((nios2_fpu_burst_6_downstream_saved_grant_ipl_memory_s1 OR nios2_fpu_burst_7_downstream_saved_grant_ipl_memory_s1) OR nios2_fpu_burst_6_downstream_saved_grant_ipl_memory_s1) OR nios2_fpu_burst_7_downstream_saved_grant_ipl_memory_s1;
  --ipl_memory_s1_arb_share_counter_next_value assignment, which is an e_assign
  ipl_memory_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(ipl_memory_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (ipl_memory_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(ipl_memory_s1_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (ipl_memory_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 4);
  --ipl_memory_s1_allgrants all slave grants, which is an e_mux
  ipl_memory_s1_allgrants <= (((or_reduce(ipl_memory_s1_grant_vector)) OR (or_reduce(ipl_memory_s1_grant_vector))) OR (or_reduce(ipl_memory_s1_grant_vector))) OR (or_reduce(ipl_memory_s1_grant_vector));
  --ipl_memory_s1_end_xfer assignment, which is an e_assign
  ipl_memory_s1_end_xfer <= NOT ((ipl_memory_s1_waits_for_read OR ipl_memory_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_ipl_memory_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_ipl_memory_s1 <= ipl_memory_s1_end_xfer AND (((NOT ipl_memory_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --ipl_memory_s1_arb_share_counter arbitration counter enable, which is an e_assign
  ipl_memory_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_ipl_memory_s1 AND ipl_memory_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_ipl_memory_s1 AND NOT ipl_memory_s1_non_bursting_master_requests));
  --ipl_memory_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ipl_memory_s1_arb_share_counter <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(ipl_memory_s1_arb_counter_enable) = '1' then 
        ipl_memory_s1_arb_share_counter <= ipl_memory_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --ipl_memory_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ipl_memory_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(ipl_memory_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_ipl_memory_s1)) OR ((end_xfer_arb_share_counter_term_ipl_memory_s1 AND NOT ipl_memory_s1_non_bursting_master_requests)))) = '1' then 
        ipl_memory_s1_slavearbiterlockenable <= or_reduce(ipl_memory_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --nios2_fpu_burst_6/downstream ipl_memory/s1 arbiterlock, which is an e_assign
  nios2_fpu_burst_6_downstream_arbiterlock <= ipl_memory_s1_slavearbiterlockenable AND nios2_fpu_burst_6_downstream_continuerequest;
  --ipl_memory_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  ipl_memory_s1_slavearbiterlockenable2 <= or_reduce(ipl_memory_s1_arb_share_counter_next_value);
  --nios2_fpu_burst_6/downstream ipl_memory/s1 arbiterlock2, which is an e_assign
  nios2_fpu_burst_6_downstream_arbiterlock2 <= ipl_memory_s1_slavearbiterlockenable2 AND nios2_fpu_burst_6_downstream_continuerequest;
  --nios2_fpu_burst_7/downstream ipl_memory/s1 arbiterlock, which is an e_assign
  nios2_fpu_burst_7_downstream_arbiterlock <= ipl_memory_s1_slavearbiterlockenable AND nios2_fpu_burst_7_downstream_continuerequest;
  --nios2_fpu_burst_7/downstream ipl_memory/s1 arbiterlock2, which is an e_assign
  nios2_fpu_burst_7_downstream_arbiterlock2 <= ipl_memory_s1_slavearbiterlockenable2 AND nios2_fpu_burst_7_downstream_continuerequest;
  --nios2_fpu_burst_7/downstream granted ipl_memory/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_nios2_fpu_burst_7_downstream_granted_slave_ipl_memory_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_nios2_fpu_burst_7_downstream_granted_slave_ipl_memory_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_7_downstream_saved_grant_ipl_memory_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ipl_memory_s1_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_7_downstream_granted_slave_ipl_memory_s1))))));
    end if;

  end process;

  --nios2_fpu_burst_7_downstream_continuerequest continued request, which is an e_mux
  nios2_fpu_burst_7_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_7_downstream_granted_slave_ipl_memory_s1))) AND std_logic_vector'("00000000000000000000000000000001")));
  --ipl_memory_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  ipl_memory_s1_any_continuerequest <= nios2_fpu_burst_7_downstream_continuerequest OR nios2_fpu_burst_6_downstream_continuerequest;
  internal_nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1 <= internal_nios2_fpu_burst_6_downstream_requests_ipl_memory_s1 AND NOT (nios2_fpu_burst_7_downstream_arbiterlock);
  --nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1_shift_register_in <= (internal_nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 AND nios2_fpu_burst_6_downstream_read) AND NOT ipl_memory_s1_waits_for_read;
  --shift register p1 nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1_shift_register) & A_ToStdLogicVector(nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1_shift_register_in)));
  --nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1_shift_register <= p1_nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1_shift_register;
    end if;

  end process;

  --local readdatavalid nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1, which is an e_mux
  nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1 <= nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1_shift_register;
  --ipl_memory_s1_writedata mux, which is an e_mux
  ipl_memory_s1_writedata <= A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_6_downstream_granted_ipl_memory_s1)) = '1'), nios2_fpu_burst_6_downstream_writedata, nios2_fpu_burst_7_downstream_writedata);
  --mux ipl_memory_s1_clken, which is an e_mux
  ipl_memory_s1_clken <= std_logic'('1');
  internal_nios2_fpu_burst_7_downstream_requests_ipl_memory_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_7_downstream_read OR nios2_fpu_burst_7_downstream_write)))))));
  --nios2_fpu_burst_6/downstream granted ipl_memory/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_nios2_fpu_burst_6_downstream_granted_slave_ipl_memory_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_nios2_fpu_burst_6_downstream_granted_slave_ipl_memory_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_6_downstream_saved_grant_ipl_memory_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ipl_memory_s1_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_6_downstream_granted_slave_ipl_memory_s1))))));
    end if;

  end process;

  --nios2_fpu_burst_6_downstream_continuerequest continued request, which is an e_mux
  nios2_fpu_burst_6_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_6_downstream_granted_slave_ipl_memory_s1))) AND std_logic_vector'("00000000000000000000000000000001")));
  internal_nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1 <= internal_nios2_fpu_burst_7_downstream_requests_ipl_memory_s1 AND NOT (nios2_fpu_burst_6_downstream_arbiterlock);
  --nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1_shift_register_in <= (internal_nios2_fpu_burst_7_downstream_granted_ipl_memory_s1 AND nios2_fpu_burst_7_downstream_read) AND NOT ipl_memory_s1_waits_for_read;
  --shift register p1 nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1_shift_register) & A_ToStdLogicVector(nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1_shift_register_in)));
  --nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1_shift_register <= p1_nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1_shift_register;
    end if;

  end process;

  --local readdatavalid nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1, which is an e_mux
  nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1 <= nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1_shift_register;
  --allow new arb cycle for ipl_memory/s1, which is an e_assign
  ipl_memory_s1_allow_new_arb_cycle <= NOT nios2_fpu_burst_6_downstream_arbiterlock AND NOT nios2_fpu_burst_7_downstream_arbiterlock;
  --nios2_fpu_burst_7/downstream assignment into master qualified-requests vector for ipl_memory/s1, which is an e_assign
  ipl_memory_s1_master_qreq_vector(0) <= internal_nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1;
  --nios2_fpu_burst_7/downstream grant ipl_memory/s1, which is an e_assign
  internal_nios2_fpu_burst_7_downstream_granted_ipl_memory_s1 <= ipl_memory_s1_grant_vector(0);
  --nios2_fpu_burst_7/downstream saved-grant ipl_memory/s1, which is an e_assign
  nios2_fpu_burst_7_downstream_saved_grant_ipl_memory_s1 <= ipl_memory_s1_arb_winner(0);
  --nios2_fpu_burst_6/downstream assignment into master qualified-requests vector for ipl_memory/s1, which is an e_assign
  ipl_memory_s1_master_qreq_vector(1) <= internal_nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1;
  --nios2_fpu_burst_6/downstream grant ipl_memory/s1, which is an e_assign
  internal_nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 <= ipl_memory_s1_grant_vector(1);
  --nios2_fpu_burst_6/downstream saved-grant ipl_memory/s1, which is an e_assign
  nios2_fpu_burst_6_downstream_saved_grant_ipl_memory_s1 <= ipl_memory_s1_arb_winner(1);
  --ipl_memory/s1 chosen-master double-vector, which is an e_assign
  ipl_memory_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((ipl_memory_s1_master_qreq_vector & ipl_memory_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT ipl_memory_s1_master_qreq_vector & NOT ipl_memory_s1_master_qreq_vector))) + (std_logic_vector'("000") & (ipl_memory_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  ipl_memory_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((ipl_memory_s1_allow_new_arb_cycle AND or_reduce(ipl_memory_s1_grant_vector)))) = '1'), ipl_memory_s1_grant_vector, ipl_memory_s1_saved_chosen_master_vector);
  --saved ipl_memory_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ipl_memory_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(ipl_memory_s1_allow_new_arb_cycle) = '1' then 
        ipl_memory_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(ipl_memory_s1_grant_vector)) = '1'), ipl_memory_s1_grant_vector, ipl_memory_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  ipl_memory_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((ipl_memory_s1_chosen_master_double_vector(1) OR ipl_memory_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((ipl_memory_s1_chosen_master_double_vector(0) OR ipl_memory_s1_chosen_master_double_vector(2)))));
  --ipl_memory/s1 chosen master rotated left, which is an e_assign
  ipl_memory_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(ipl_memory_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(ipl_memory_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --ipl_memory/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ipl_memory_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(ipl_memory_s1_grant_vector)) = '1' then 
        ipl_memory_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(ipl_memory_s1_end_xfer) = '1'), ipl_memory_s1_chosen_master_rot_left, ipl_memory_s1_grant_vector);
      end if;
    end if;

  end process;

  --~ipl_memory_s1_reset assignment, which is an e_assign
  ipl_memory_s1_reset <= NOT reset_n;
  ipl_memory_s1_chipselect <= internal_nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 OR internal_nios2_fpu_burst_7_downstream_granted_ipl_memory_s1;
  --ipl_memory_s1_firsttransfer first transaction, which is an e_assign
  ipl_memory_s1_firsttransfer <= A_WE_StdLogic((std_logic'(ipl_memory_s1_begins_xfer) = '1'), ipl_memory_s1_unreg_firsttransfer, ipl_memory_s1_reg_firsttransfer);
  --ipl_memory_s1_unreg_firsttransfer first transaction, which is an e_assign
  ipl_memory_s1_unreg_firsttransfer <= NOT ((ipl_memory_s1_slavearbiterlockenable AND ipl_memory_s1_any_continuerequest));
  --ipl_memory_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ipl_memory_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(ipl_memory_s1_begins_xfer) = '1' then 
        ipl_memory_s1_reg_firsttransfer <= ipl_memory_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --ipl_memory_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  ipl_memory_s1_beginbursttransfer_internal <= ipl_memory_s1_begins_xfer;
  --ipl_memory_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  ipl_memory_s1_arbitration_holdoff_internal <= ipl_memory_s1_begins_xfer AND ipl_memory_s1_firsttransfer;
  --ipl_memory_s1_write assignment, which is an e_mux
  ipl_memory_s1_write <= ((internal_nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 AND nios2_fpu_burst_6_downstream_write)) OR ((internal_nios2_fpu_burst_7_downstream_granted_ipl_memory_s1 AND nios2_fpu_burst_7_downstream_write));
  shifted_address_to_ipl_memory_s1_from_nios2_fpu_burst_6_downstream <= nios2_fpu_burst_6_downstream_address_to_slave;
  --ipl_memory_s1_address mux, which is an e_mux
  ipl_memory_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_6_downstream_granted_ipl_memory_s1)) = '1'), (A_SRL(shifted_address_to_ipl_memory_s1_from_nios2_fpu_burst_6_downstream,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_ipl_memory_s1_from_nios2_fpu_burst_7_downstream,std_logic_vector'("00000000000000000000000000000010")))), 11);
  shifted_address_to_ipl_memory_s1_from_nios2_fpu_burst_7_downstream <= nios2_fpu_burst_7_downstream_address_to_slave;
  --d1_ipl_memory_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_ipl_memory_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_ipl_memory_s1_end_xfer <= ipl_memory_s1_end_xfer;
    end if;

  end process;

  --ipl_memory_s1_waits_for_read in a cycle, which is an e_mux
  ipl_memory_s1_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ipl_memory_s1_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --ipl_memory_s1_in_a_read_cycle assignment, which is an e_assign
  ipl_memory_s1_in_a_read_cycle <= ((internal_nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 AND nios2_fpu_burst_6_downstream_read)) OR ((internal_nios2_fpu_burst_7_downstream_granted_ipl_memory_s1 AND nios2_fpu_burst_7_downstream_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= ipl_memory_s1_in_a_read_cycle;
  --ipl_memory_s1_waits_for_write in a cycle, which is an e_mux
  ipl_memory_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ipl_memory_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --ipl_memory_s1_in_a_write_cycle assignment, which is an e_assign
  ipl_memory_s1_in_a_write_cycle <= ((internal_nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 AND nios2_fpu_burst_6_downstream_write)) OR ((internal_nios2_fpu_burst_7_downstream_granted_ipl_memory_s1 AND nios2_fpu_burst_7_downstream_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= ipl_memory_s1_in_a_write_cycle;
  wait_for_ipl_memory_s1_counter <= std_logic'('0');
  --ipl_memory_s1_byteenable byte enable port mux, which is an e_mux
  ipl_memory_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_6_downstream_granted_ipl_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_6_downstream_byteenable)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_7_downstream_granted_ipl_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_7_downstream_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))), 4);
  --vhdl renameroo for output signals
  nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 <= internal_nios2_fpu_burst_6_downstream_granted_ipl_memory_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1 <= internal_nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_6_downstream_requests_ipl_memory_s1 <= internal_nios2_fpu_burst_6_downstream_requests_ipl_memory_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_7_downstream_granted_ipl_memory_s1 <= internal_nios2_fpu_burst_7_downstream_granted_ipl_memory_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1 <= internal_nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_7_downstream_requests_ipl_memory_s1 <= internal_nios2_fpu_burst_7_downstream_requests_ipl_memory_s1;
--synthesis translate_off
    --ipl_memory/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --nios2_fpu_burst_6/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line2 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_6_downstream_requests_ipl_memory_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_6_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line2, now);
          write(write_line2, string'(": "));
          write(write_line2, string'("nios2_fpu_burst_6/downstream drove 0 on its 'arbitrationshare' port while accessing slave ipl_memory/s1"));
          write(output, write_line2.all);
          deallocate (write_line2);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_6/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line3 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_6_downstream_requests_ipl_memory_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_6_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line3, now);
          write(write_line3, string'(": "));
          write(write_line3, string'("nios2_fpu_burst_6/downstream drove 0 on its 'burstcount' port while accessing slave ipl_memory/s1"));
          write(output, write_line3.all);
          deallocate (write_line3);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_7/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line4 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_7_downstream_requests_ipl_memory_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_7_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line4, now);
          write(write_line4, string'(": "));
          write(write_line4, string'("nios2_fpu_burst_7/downstream drove 0 on its 'arbitrationshare' port while accessing slave ipl_memory/s1"));
          write(output, write_line4.all);
          deallocate (write_line4);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_7/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line5 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_7_downstream_requests_ipl_memory_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_7_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line5, now);
          write(write_line5, string'(": "));
          write(write_line5, string'("nios2_fpu_burst_7/downstream drove 0 on its 'burstcount' port while accessing slave ipl_memory/s1"));
          write(output, write_line5.all);
          deallocate (write_line5);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line6 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_6_downstream_granted_ipl_memory_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_7_downstream_granted_ipl_memory_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line6, now);
          write(write_line6, string'(": "));
          write(write_line6, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line6.all);
          deallocate (write_line6);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line7 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_6_downstream_saved_grant_ipl_memory_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_7_downstream_saved_grant_ipl_memory_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line7, now);
          write(write_line7, string'(": "));
          write(write_line7, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line7.all);
          deallocate (write_line7);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity jtag_uart_avalon_jtag_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                 signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                 signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                 signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read : IN STD_LOGIC;
                 signal peripheral_bridge_m1_write : IN STD_LOGIC;
                 signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_jtag_uart_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_address : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC
              );
end entity jtag_uart_avalon_jtag_slave_arbitrator;


architecture europa of jtag_uart_avalon_jtag_slave_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_allgrants :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_any_continuerequest :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_counter_enable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_share_counter :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_share_set_values :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_begins_xfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_grant_vector :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_in_a_read_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_in_a_write_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_master_qreq_vector :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_non_bursting_master_requests :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_reg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_slavearbiterlockenable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_unreg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waits_for_read :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waits_for_write :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal peripheral_bridge_m1_continuerequest :  STD_LOGIC;
                signal peripheral_bridge_m1_saved_grant_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal shifted_address_to_jtag_uart_avalon_jtag_slave_from_peripheral_bridge_m1 :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal wait_for_jtag_uart_avalon_jtag_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT jtag_uart_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  jtag_uart_avalon_jtag_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave);
  --assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_readdata_from_sa <= jtag_uart_avalon_jtag_slave_readdata;
  internal_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave <= to_std_logic(((Std_Logic_Vector'(peripheral_bridge_m1_address_to_slave(12 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("0000010000000")))) AND peripheral_bridge_m1_chipselect;
  --assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_dataavailable_from_sa <= jtag_uart_avalon_jtag_slave_dataavailable;
  --assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_readyfordata_from_sa <= jtag_uart_avalon_jtag_slave_readyfordata;
  --assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa <= jtag_uart_avalon_jtag_slave_waitrequest;
  --jtag_uart_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  jtag_uart_avalon_jtag_slave_arb_share_set_values <= std_logic'('1');
  --jtag_uart_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_non_bursting_master_requests <= internal_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  --jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --jtag_uart_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(jtag_uart_avalon_jtag_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(jtag_uart_avalon_jtag_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(jtag_uart_avalon_jtag_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(jtag_uart_avalon_jtag_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --jtag_uart_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  jtag_uart_avalon_jtag_slave_allgrants <= jtag_uart_avalon_jtag_slave_grant_vector;
  --jtag_uart_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_end_xfer <= NOT ((jtag_uart_avalon_jtag_slave_waits_for_read OR jtag_uart_avalon_jtag_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave <= jtag_uart_avalon_jtag_slave_end_xfer AND (((NOT jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --jtag_uart_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  jtag_uart_avalon_jtag_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND jtag_uart_avalon_jtag_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND NOT jtag_uart_avalon_jtag_slave_non_bursting_master_requests));
  --jtag_uart_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_avalon_jtag_slave_arb_counter_enable) = '1' then 
        jtag_uart_avalon_jtag_slave_arb_share_counter <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((jtag_uart_avalon_jtag_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave)) OR ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND NOT jtag_uart_avalon_jtag_slave_non_bursting_master_requests)))) = '1' then 
        jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --peripheral_bridge/m1 jtag_uart/avalon_jtag_slave arbiterlock, which is an e_assign
  peripheral_bridge_m1_arbiterlock <= jtag_uart_avalon_jtag_slave_slavearbiterlockenable AND peripheral_bridge_m1_continuerequest;
  --jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
  --peripheral_bridge/m1 jtag_uart/avalon_jtag_slave arbiterlock2, which is an e_assign
  peripheral_bridge_m1_arbiterlock2 <= jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 AND peripheral_bridge_m1_continuerequest;
  --jtag_uart_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  jtag_uart_avalon_jtag_slave_any_continuerequest <= std_logic'('1');
  --peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  peripheral_bridge_m1_continuerequest <= std_logic'('1');
  internal_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave <= internal_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave AND NOT ((((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave, which is an e_mux
  peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave <= (internal_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect))) AND NOT jtag_uart_avalon_jtag_slave_waits_for_read;
  --jtag_uart_avalon_jtag_slave_writedata mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_writedata <= peripheral_bridge_m1_writedata;
  --master is always granted when requested
  internal_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave <= internal_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  --peripheral_bridge/m1 saved-grant jtag_uart/avalon_jtag_slave, which is an e_assign
  peripheral_bridge_m1_saved_grant_jtag_uart_avalon_jtag_slave <= internal_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  --allow new arb cycle for jtag_uart/avalon_jtag_slave, which is an e_assign
  jtag_uart_avalon_jtag_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  jtag_uart_avalon_jtag_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  jtag_uart_avalon_jtag_slave_master_qreq_vector <= std_logic'('1');
  --jtag_uart_avalon_jtag_slave_reset_n assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_reset_n <= reset_n;
  jtag_uart_avalon_jtag_slave_chipselect <= internal_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  --jtag_uart_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  jtag_uart_avalon_jtag_slave_firsttransfer <= A_WE_StdLogic((std_logic'(jtag_uart_avalon_jtag_slave_begins_xfer) = '1'), jtag_uart_avalon_jtag_slave_unreg_firsttransfer, jtag_uart_avalon_jtag_slave_reg_firsttransfer);
  --jtag_uart_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  jtag_uart_avalon_jtag_slave_unreg_firsttransfer <= NOT ((jtag_uart_avalon_jtag_slave_slavearbiterlockenable AND jtag_uart_avalon_jtag_slave_any_continuerequest));
  --jtag_uart_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_avalon_jtag_slave_begins_xfer) = '1' then 
        jtag_uart_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  jtag_uart_avalon_jtag_slave_beginbursttransfer_internal <= jtag_uart_avalon_jtag_slave_begins_xfer;
  --~jtag_uart_avalon_jtag_slave_read_n assignment, which is an e_mux
  jtag_uart_avalon_jtag_slave_read_n <= NOT ((internal_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect))));
  --~jtag_uart_avalon_jtag_slave_write_n assignment, which is an e_mux
  jtag_uart_avalon_jtag_slave_write_n <= NOT ((internal_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect))));
  shifted_address_to_jtag_uart_avalon_jtag_slave_from_peripheral_bridge_m1 <= peripheral_bridge_m1_address_to_slave;
  --jtag_uart_avalon_jtag_slave_address mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_address <= Vector_To_Std_Logic(A_SRL(shifted_address_to_jtag_uart_avalon_jtag_slave_from_peripheral_bridge_m1,std_logic_vector'("00000000000000000000000000000010")));
  --d1_jtag_uart_avalon_jtag_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_jtag_uart_avalon_jtag_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_jtag_uart_avalon_jtag_slave_end_xfer <= jtag_uart_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  jtag_uart_avalon_jtag_slave_waits_for_read <= jtag_uart_avalon_jtag_slave_in_a_read_cycle AND internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_in_a_read_cycle <= internal_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= jtag_uart_avalon_jtag_slave_in_a_read_cycle;
  --jtag_uart_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  jtag_uart_avalon_jtag_slave_waits_for_write <= jtag_uart_avalon_jtag_slave_in_a_write_cycle AND internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_in_a_write_cycle <= internal_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= jtag_uart_avalon_jtag_slave_in_a_write_cycle;
  wait_for_jtag_uart_avalon_jtag_slave_counter <= std_logic'('0');
  --assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_irq_from_sa <= jtag_uart_avalon_jtag_slave_irq;
  --vhdl renameroo for output signals
  jtag_uart_avalon_jtag_slave_waitrequest_from_sa <= internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave <= internal_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave <= internal_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave <= internal_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
--synthesis translate_off
    --jtag_uart/avalon_jtag_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --peripheral_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line8 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line8, now);
          write(write_line8, string'(": "));
          write(write_line8, string'("peripheral_bridge/m1 drove 0 on its 'burstcount' port while accessing slave jtag_uart/avalon_jtag_slave"));
          write(output, write_line8.all);
          deallocate (write_line8);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity led_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal led_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                 signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                 signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read : IN STD_LOGIC;
                 signal peripheral_bridge_m1_write : IN STD_LOGIC;
                 signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_led_s1_end_xfer : OUT STD_LOGIC;
                 signal led_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal led_s1_chipselect : OUT STD_LOGIC;
                 signal led_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal led_s1_reset_n : OUT STD_LOGIC;
                 signal led_s1_write_n : OUT STD_LOGIC;
                 signal led_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal peripheral_bridge_m1_granted_led_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_led_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_led_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_requests_led_s1 : OUT STD_LOGIC
              );
end entity led_s1_arbitrator;


architecture europa of led_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_led_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_granted_led_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_qualified_request_led_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_requests_led_s1 :  STD_LOGIC;
                signal led_s1_allgrants :  STD_LOGIC;
                signal led_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal led_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal led_s1_any_continuerequest :  STD_LOGIC;
                signal led_s1_arb_counter_enable :  STD_LOGIC;
                signal led_s1_arb_share_counter :  STD_LOGIC;
                signal led_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal led_s1_arb_share_set_values :  STD_LOGIC;
                signal led_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal led_s1_begins_xfer :  STD_LOGIC;
                signal led_s1_end_xfer :  STD_LOGIC;
                signal led_s1_firsttransfer :  STD_LOGIC;
                signal led_s1_grant_vector :  STD_LOGIC;
                signal led_s1_in_a_read_cycle :  STD_LOGIC;
                signal led_s1_in_a_write_cycle :  STD_LOGIC;
                signal led_s1_master_qreq_vector :  STD_LOGIC;
                signal led_s1_non_bursting_master_requests :  STD_LOGIC;
                signal led_s1_reg_firsttransfer :  STD_LOGIC;
                signal led_s1_slavearbiterlockenable :  STD_LOGIC;
                signal led_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal led_s1_unreg_firsttransfer :  STD_LOGIC;
                signal led_s1_waits_for_read :  STD_LOGIC;
                signal led_s1_waits_for_write :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal peripheral_bridge_m1_continuerequest :  STD_LOGIC;
                signal peripheral_bridge_m1_saved_grant_led_s1 :  STD_LOGIC;
                signal shifted_address_to_led_s1_from_peripheral_bridge_m1 :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal wait_for_led_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT led_s1_end_xfer;
    end if;

  end process;

  led_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_peripheral_bridge_m1_qualified_request_led_s1);
  --assign led_s1_readdata_from_sa = led_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  led_s1_readdata_from_sa <= led_s1_readdata;
  internal_peripheral_bridge_m1_requests_led_s1 <= to_std_logic(((Std_Logic_Vector'(peripheral_bridge_m1_address_to_slave(12 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("0001000000000")))) AND peripheral_bridge_m1_chipselect;
  --led_s1_arb_share_counter set values, which is an e_mux
  led_s1_arb_share_set_values <= std_logic'('1');
  --led_s1_non_bursting_master_requests mux, which is an e_mux
  led_s1_non_bursting_master_requests <= internal_peripheral_bridge_m1_requests_led_s1;
  --led_s1_any_bursting_master_saved_grant mux, which is an e_mux
  led_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --led_s1_arb_share_counter_next_value assignment, which is an e_assign
  led_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(led_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(led_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(led_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(led_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --led_s1_allgrants all slave grants, which is an e_mux
  led_s1_allgrants <= led_s1_grant_vector;
  --led_s1_end_xfer assignment, which is an e_assign
  led_s1_end_xfer <= NOT ((led_s1_waits_for_read OR led_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_led_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_led_s1 <= led_s1_end_xfer AND (((NOT led_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --led_s1_arb_share_counter arbitration counter enable, which is an e_assign
  led_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_led_s1 AND led_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_led_s1 AND NOT led_s1_non_bursting_master_requests));
  --led_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      led_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(led_s1_arb_counter_enable) = '1' then 
        led_s1_arb_share_counter <= led_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --led_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      led_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((led_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_led_s1)) OR ((end_xfer_arb_share_counter_term_led_s1 AND NOT led_s1_non_bursting_master_requests)))) = '1' then 
        led_s1_slavearbiterlockenable <= led_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --peripheral_bridge/m1 led/s1 arbiterlock, which is an e_assign
  peripheral_bridge_m1_arbiterlock <= led_s1_slavearbiterlockenable AND peripheral_bridge_m1_continuerequest;
  --led_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  led_s1_slavearbiterlockenable2 <= led_s1_arb_share_counter_next_value;
  --peripheral_bridge/m1 led/s1 arbiterlock2, which is an e_assign
  peripheral_bridge_m1_arbiterlock2 <= led_s1_slavearbiterlockenable2 AND peripheral_bridge_m1_continuerequest;
  --led_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  led_s1_any_continuerequest <= std_logic'('1');
  --peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  peripheral_bridge_m1_continuerequest <= std_logic'('1');
  internal_peripheral_bridge_m1_qualified_request_led_s1 <= internal_peripheral_bridge_m1_requests_led_s1 AND NOT ((((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid peripheral_bridge_m1_read_data_valid_led_s1, which is an e_mux
  peripheral_bridge_m1_read_data_valid_led_s1 <= (internal_peripheral_bridge_m1_granted_led_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect))) AND NOT led_s1_waits_for_read;
  --led_s1_writedata mux, which is an e_mux
  led_s1_writedata <= peripheral_bridge_m1_writedata;
  --master is always granted when requested
  internal_peripheral_bridge_m1_granted_led_s1 <= internal_peripheral_bridge_m1_qualified_request_led_s1;
  --peripheral_bridge/m1 saved-grant led/s1, which is an e_assign
  peripheral_bridge_m1_saved_grant_led_s1 <= internal_peripheral_bridge_m1_requests_led_s1;
  --allow new arb cycle for led/s1, which is an e_assign
  led_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  led_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  led_s1_master_qreq_vector <= std_logic'('1');
  --led_s1_reset_n assignment, which is an e_assign
  led_s1_reset_n <= reset_n;
  led_s1_chipselect <= internal_peripheral_bridge_m1_granted_led_s1;
  --led_s1_firsttransfer first transaction, which is an e_assign
  led_s1_firsttransfer <= A_WE_StdLogic((std_logic'(led_s1_begins_xfer) = '1'), led_s1_unreg_firsttransfer, led_s1_reg_firsttransfer);
  --led_s1_unreg_firsttransfer first transaction, which is an e_assign
  led_s1_unreg_firsttransfer <= NOT ((led_s1_slavearbiterlockenable AND led_s1_any_continuerequest));
  --led_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      led_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(led_s1_begins_xfer) = '1' then 
        led_s1_reg_firsttransfer <= led_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --led_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  led_s1_beginbursttransfer_internal <= led_s1_begins_xfer;
  --~led_s1_write_n assignment, which is an e_mux
  led_s1_write_n <= NOT ((internal_peripheral_bridge_m1_granted_led_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect))));
  shifted_address_to_led_s1_from_peripheral_bridge_m1 <= peripheral_bridge_m1_address_to_slave;
  --led_s1_address mux, which is an e_mux
  led_s1_address <= A_EXT (A_SRL(shifted_address_to_led_s1_from_peripheral_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_led_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_led_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_led_s1_end_xfer <= led_s1_end_xfer;
    end if;

  end process;

  --led_s1_waits_for_read in a cycle, which is an e_mux
  led_s1_waits_for_read <= led_s1_in_a_read_cycle AND led_s1_begins_xfer;
  --led_s1_in_a_read_cycle assignment, which is an e_assign
  led_s1_in_a_read_cycle <= internal_peripheral_bridge_m1_granted_led_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= led_s1_in_a_read_cycle;
  --led_s1_waits_for_write in a cycle, which is an e_mux
  led_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(led_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --led_s1_in_a_write_cycle assignment, which is an e_assign
  led_s1_in_a_write_cycle <= internal_peripheral_bridge_m1_granted_led_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= led_s1_in_a_write_cycle;
  wait_for_led_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  peripheral_bridge_m1_granted_led_s1 <= internal_peripheral_bridge_m1_granted_led_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_qualified_request_led_s1 <= internal_peripheral_bridge_m1_qualified_request_led_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_requests_led_s1 <= internal_peripheral_bridge_m1_requests_led_s1;
--synthesis translate_off
    --led/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --peripheral_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line9 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_peripheral_bridge_m1_requests_led_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line9, now);
          write(write_line9, string'(": "));
          write(write_line9, string'("peripheral_bridge/m1 drove 0 on its 'burstcount' port while accessing slave led/s1"));
          write(output, write_line9.all);
          deallocate (write_line9);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity mmcdma_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal mmcdma_s1_irq : IN STD_LOGIC;
                 signal mmcdma_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                 signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                 signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read : IN STD_LOGIC;
                 signal peripheral_bridge_m1_write : IN STD_LOGIC;
                 signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_mmcdma_s1_end_xfer : OUT STD_LOGIC;
                 signal mmcdma_s1_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal mmcdma_s1_chipselect : OUT STD_LOGIC;
                 signal mmcdma_s1_irq_from_sa : OUT STD_LOGIC;
                 signal mmcdma_s1_read : OUT STD_LOGIC;
                 signal mmcdma_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal mmcdma_s1_reset : OUT STD_LOGIC;
                 signal mmcdma_s1_wait_counter_eq_0 : OUT STD_LOGIC;
                 signal mmcdma_s1_write : OUT STD_LOGIC;
                 signal mmcdma_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal peripheral_bridge_m1_granted_mmcdma_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_mmcdma_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_mmcdma_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_requests_mmcdma_s1 : OUT STD_LOGIC
              );
end entity mmcdma_s1_arbitrator;


architecture europa of mmcdma_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_mmcdma_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_mmcdma_s1_wait_counter_eq_0 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_granted_mmcdma_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_qualified_request_mmcdma_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_requests_mmcdma_s1 :  STD_LOGIC;
                signal mmcdma_s1_allgrants :  STD_LOGIC;
                signal mmcdma_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal mmcdma_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal mmcdma_s1_any_continuerequest :  STD_LOGIC;
                signal mmcdma_s1_arb_counter_enable :  STD_LOGIC;
                signal mmcdma_s1_arb_share_counter :  STD_LOGIC;
                signal mmcdma_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal mmcdma_s1_arb_share_set_values :  STD_LOGIC;
                signal mmcdma_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal mmcdma_s1_begins_xfer :  STD_LOGIC;
                signal mmcdma_s1_counter_load_value :  STD_LOGIC;
                signal mmcdma_s1_end_xfer :  STD_LOGIC;
                signal mmcdma_s1_firsttransfer :  STD_LOGIC;
                signal mmcdma_s1_grant_vector :  STD_LOGIC;
                signal mmcdma_s1_in_a_read_cycle :  STD_LOGIC;
                signal mmcdma_s1_in_a_write_cycle :  STD_LOGIC;
                signal mmcdma_s1_master_qreq_vector :  STD_LOGIC;
                signal mmcdma_s1_non_bursting_master_requests :  STD_LOGIC;
                signal mmcdma_s1_reg_firsttransfer :  STD_LOGIC;
                signal mmcdma_s1_slavearbiterlockenable :  STD_LOGIC;
                signal mmcdma_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal mmcdma_s1_unreg_firsttransfer :  STD_LOGIC;
                signal mmcdma_s1_wait_counter :  STD_LOGIC;
                signal mmcdma_s1_waits_for_read :  STD_LOGIC;
                signal mmcdma_s1_waits_for_write :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal peripheral_bridge_m1_continuerequest :  STD_LOGIC;
                signal peripheral_bridge_m1_saved_grant_mmcdma_s1 :  STD_LOGIC;
                signal shifted_address_to_mmcdma_s1_from_peripheral_bridge_m1 :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal wait_for_mmcdma_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT mmcdma_s1_end_xfer;
    end if;

  end process;

  mmcdma_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_peripheral_bridge_m1_qualified_request_mmcdma_s1);
  --assign mmcdma_s1_readdata_from_sa = mmcdma_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  mmcdma_s1_readdata_from_sa <= mmcdma_s1_readdata;
  internal_peripheral_bridge_m1_requests_mmcdma_s1 <= to_std_logic(((Std_Logic_Vector'(peripheral_bridge_m1_address_to_slave(12 DOWNTO 10) & std_logic_vector'("0000000000")) = std_logic_vector'("0010000000000")))) AND peripheral_bridge_m1_chipselect;
  --mmcdma_s1_arb_share_counter set values, which is an e_mux
  mmcdma_s1_arb_share_set_values <= std_logic'('1');
  --mmcdma_s1_non_bursting_master_requests mux, which is an e_mux
  mmcdma_s1_non_bursting_master_requests <= internal_peripheral_bridge_m1_requests_mmcdma_s1;
  --mmcdma_s1_any_bursting_master_saved_grant mux, which is an e_mux
  mmcdma_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --mmcdma_s1_arb_share_counter_next_value assignment, which is an e_assign
  mmcdma_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(mmcdma_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(mmcdma_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(mmcdma_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(mmcdma_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --mmcdma_s1_allgrants all slave grants, which is an e_mux
  mmcdma_s1_allgrants <= mmcdma_s1_grant_vector;
  --mmcdma_s1_end_xfer assignment, which is an e_assign
  mmcdma_s1_end_xfer <= NOT ((mmcdma_s1_waits_for_read OR mmcdma_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_mmcdma_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_mmcdma_s1 <= mmcdma_s1_end_xfer AND (((NOT mmcdma_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --mmcdma_s1_arb_share_counter arbitration counter enable, which is an e_assign
  mmcdma_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_mmcdma_s1 AND mmcdma_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_mmcdma_s1 AND NOT mmcdma_s1_non_bursting_master_requests));
  --mmcdma_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      mmcdma_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(mmcdma_s1_arb_counter_enable) = '1' then 
        mmcdma_s1_arb_share_counter <= mmcdma_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --mmcdma_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      mmcdma_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((mmcdma_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_mmcdma_s1)) OR ((end_xfer_arb_share_counter_term_mmcdma_s1 AND NOT mmcdma_s1_non_bursting_master_requests)))) = '1' then 
        mmcdma_s1_slavearbiterlockenable <= mmcdma_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --peripheral_bridge/m1 mmcdma/s1 arbiterlock, which is an e_assign
  peripheral_bridge_m1_arbiterlock <= mmcdma_s1_slavearbiterlockenable AND peripheral_bridge_m1_continuerequest;
  --mmcdma_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  mmcdma_s1_slavearbiterlockenable2 <= mmcdma_s1_arb_share_counter_next_value;
  --peripheral_bridge/m1 mmcdma/s1 arbiterlock2, which is an e_assign
  peripheral_bridge_m1_arbiterlock2 <= mmcdma_s1_slavearbiterlockenable2 AND peripheral_bridge_m1_continuerequest;
  --mmcdma_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  mmcdma_s1_any_continuerequest <= std_logic'('1');
  --peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  peripheral_bridge_m1_continuerequest <= std_logic'('1');
  internal_peripheral_bridge_m1_qualified_request_mmcdma_s1 <= internal_peripheral_bridge_m1_requests_mmcdma_s1 AND NOT ((((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid peripheral_bridge_m1_read_data_valid_mmcdma_s1, which is an e_mux
  peripheral_bridge_m1_read_data_valid_mmcdma_s1 <= (internal_peripheral_bridge_m1_granted_mmcdma_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect))) AND NOT mmcdma_s1_waits_for_read;
  --mmcdma_s1_writedata mux, which is an e_mux
  mmcdma_s1_writedata <= peripheral_bridge_m1_writedata;
  --master is always granted when requested
  internal_peripheral_bridge_m1_granted_mmcdma_s1 <= internal_peripheral_bridge_m1_qualified_request_mmcdma_s1;
  --peripheral_bridge/m1 saved-grant mmcdma/s1, which is an e_assign
  peripheral_bridge_m1_saved_grant_mmcdma_s1 <= internal_peripheral_bridge_m1_requests_mmcdma_s1;
  --allow new arb cycle for mmcdma/s1, which is an e_assign
  mmcdma_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  mmcdma_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  mmcdma_s1_master_qreq_vector <= std_logic'('1');
  --~mmcdma_s1_reset assignment, which is an e_assign
  mmcdma_s1_reset <= NOT reset_n;
  mmcdma_s1_chipselect <= internal_peripheral_bridge_m1_granted_mmcdma_s1;
  --mmcdma_s1_firsttransfer first transaction, which is an e_assign
  mmcdma_s1_firsttransfer <= A_WE_StdLogic((std_logic'(mmcdma_s1_begins_xfer) = '1'), mmcdma_s1_unreg_firsttransfer, mmcdma_s1_reg_firsttransfer);
  --mmcdma_s1_unreg_firsttransfer first transaction, which is an e_assign
  mmcdma_s1_unreg_firsttransfer <= NOT ((mmcdma_s1_slavearbiterlockenable AND mmcdma_s1_any_continuerequest));
  --mmcdma_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      mmcdma_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(mmcdma_s1_begins_xfer) = '1' then 
        mmcdma_s1_reg_firsttransfer <= mmcdma_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --mmcdma_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  mmcdma_s1_beginbursttransfer_internal <= mmcdma_s1_begins_xfer;
  --mmcdma_s1_read assignment, which is an e_mux
  mmcdma_s1_read <= internal_peripheral_bridge_m1_granted_mmcdma_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --mmcdma_s1_write assignment, which is an e_mux
  mmcdma_s1_write <= internal_peripheral_bridge_m1_granted_mmcdma_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect));
  shifted_address_to_mmcdma_s1_from_peripheral_bridge_m1 <= peripheral_bridge_m1_address_to_slave;
  --mmcdma_s1_address mux, which is an e_mux
  mmcdma_s1_address <= A_EXT (A_SRL(shifted_address_to_mmcdma_s1_from_peripheral_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 8);
  --d1_mmcdma_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_mmcdma_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_mmcdma_s1_end_xfer <= mmcdma_s1_end_xfer;
    end if;

  end process;

  --mmcdma_s1_waits_for_read in a cycle, which is an e_mux
  mmcdma_s1_waits_for_read <= mmcdma_s1_in_a_read_cycle AND wait_for_mmcdma_s1_counter;
  --mmcdma_s1_in_a_read_cycle assignment, which is an e_assign
  mmcdma_s1_in_a_read_cycle <= internal_peripheral_bridge_m1_granted_mmcdma_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= mmcdma_s1_in_a_read_cycle;
  --mmcdma_s1_waits_for_write in a cycle, which is an e_mux
  mmcdma_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(mmcdma_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --mmcdma_s1_in_a_write_cycle assignment, which is an e_assign
  mmcdma_s1_in_a_write_cycle <= internal_peripheral_bridge_m1_granted_mmcdma_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= mmcdma_s1_in_a_write_cycle;
  internal_mmcdma_s1_wait_counter_eq_0 <= to_std_logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(mmcdma_s1_wait_counter))) = std_logic_vector'("00000000000000000000000000000000")));
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      mmcdma_s1_wait_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      mmcdma_s1_wait_counter <= mmcdma_s1_counter_load_value;
    end if;

  end process;

  mmcdma_s1_counter_load_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((mmcdma_s1_in_a_read_cycle AND mmcdma_s1_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'((NOT internal_mmcdma_s1_wait_counter_eq_0)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(mmcdma_s1_wait_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  wait_for_mmcdma_s1_counter <= mmcdma_s1_begins_xfer OR NOT internal_mmcdma_s1_wait_counter_eq_0;
  --assign mmcdma_s1_irq_from_sa = mmcdma_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  mmcdma_s1_irq_from_sa <= mmcdma_s1_irq;
  --vhdl renameroo for output signals
  mmcdma_s1_wait_counter_eq_0 <= internal_mmcdma_s1_wait_counter_eq_0;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_granted_mmcdma_s1 <= internal_peripheral_bridge_m1_granted_mmcdma_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_qualified_request_mmcdma_s1 <= internal_peripheral_bridge_m1_qualified_request_mmcdma_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_requests_mmcdma_s1 <= internal_peripheral_bridge_m1_requests_mmcdma_s1;
--synthesis translate_off
    --mmcdma/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --peripheral_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line10 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_peripheral_bridge_m1_requests_mmcdma_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line10, now);
          write(write_line10, string'(": "));
          write(write_line10, string'("peripheral_bridge/m1 drove 0 on its 'burstcount' port while accessing slave mmcdma/s1"));
          write(output, write_line10.all);
          deallocate (write_line10);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fast_fpu_jtag_debug_module_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fast_fpu_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_jtag_debug_module_resetrequest : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_address_to_slave : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal nios2_fpu_burst_4_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_4_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_4_downstream_debugaccess : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_latency_counter : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_5_downstream_address_to_slave : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal nios2_fpu_burst_5_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_5_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_5_downstream_debugaccess : IN STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_latency_counter : IN STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_nios2_fast_fpu_jtag_debug_module_end_xfer : OUT STD_LOGIC;
                 signal nios2_fast_fpu_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                 signal nios2_fast_fpu_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                 signal nios2_fast_fpu_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fast_fpu_jtag_debug_module_chipselect : OUT STD_LOGIC;
                 signal nios2_fast_fpu_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                 signal nios2_fast_fpu_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_fast_fpu_jtag_debug_module_write : OUT STD_LOGIC;
                 signal nios2_fast_fpu_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC
              );
end entity nios2_fast_fpu_jtag_debug_module_arbitrator;


architecture europa of nios2_fast_fpu_jtag_debug_module_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal internal_nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal internal_nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal internal_nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal internal_nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal internal_nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_nios2_fpu_burst_4_downstream_granted_slave_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_nios2_fpu_burst_5_downstream_granted_slave_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_allgrants :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_any_continuerequest :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_jtag_debug_module_arb_counter_enable :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_arb_share_counter :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fast_fpu_jtag_debug_module_arb_share_counter_next_value :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fast_fpu_jtag_debug_module_arb_share_set_values :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fast_fpu_jtag_debug_module_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_jtag_debug_module_arbitration_holdoff_internal :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_begins_xfer :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fast_fpu_jtag_debug_module_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_firsttransfer :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_jtag_debug_module_in_a_read_cycle :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_in_a_write_cycle :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_jtag_debug_module_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_reg_firsttransfer :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_jtag_debug_module_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_waits_for_read :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_waits_for_write :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_arbiterlock :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_arbiterlock2 :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_saved_grant_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_arbiterlock :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_arbiterlock2 :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_saved_grant_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal shifted_address_to_nios2_fast_fpu_jtag_debug_module_from_nios2_fpu_burst_4_downstream :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal shifted_address_to_nios2_fast_fpu_jtag_debug_module_from_nios2_fpu_burst_5_downstream :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal wait_for_nios2_fast_fpu_jtag_debug_module_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_fast_fpu_jtag_debug_module_end_xfer;
    end if;

  end process;

  nios2_fast_fpu_jtag_debug_module_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module OR internal_nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module));
  --assign nios2_fast_fpu_jtag_debug_module_readdata_from_sa = nios2_fast_fpu_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_readdata_from_sa <= nios2_fast_fpu_jtag_debug_module_readdata;
  internal_nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_4_downstream_read OR nios2_fpu_burst_4_downstream_write)))))));
  --nios2_fast_fpu_jtag_debug_module_arb_share_counter set values, which is an e_mux
  nios2_fast_fpu_jtag_debug_module_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_4_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_5_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_4_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_5_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001"))))), 4);
  --nios2_fast_fpu_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  nios2_fast_fpu_jtag_debug_module_non_bursting_master_requests <= std_logic'('0');
  --nios2_fast_fpu_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_fast_fpu_jtag_debug_module_any_bursting_master_saved_grant <= ((nios2_fpu_burst_4_downstream_saved_grant_nios2_fast_fpu_jtag_debug_module OR nios2_fpu_burst_5_downstream_saved_grant_nios2_fast_fpu_jtag_debug_module) OR nios2_fpu_burst_4_downstream_saved_grant_nios2_fast_fpu_jtag_debug_module) OR nios2_fpu_burst_5_downstream_saved_grant_nios2_fast_fpu_jtag_debug_module;
  --nios2_fast_fpu_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_fast_fpu_jtag_debug_module_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (nios2_fast_fpu_jtag_debug_module_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_fast_fpu_jtag_debug_module_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (nios2_fast_fpu_jtag_debug_module_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 4);
  --nios2_fast_fpu_jtag_debug_module_allgrants all slave grants, which is an e_mux
  nios2_fast_fpu_jtag_debug_module_allgrants <= (((or_reduce(nios2_fast_fpu_jtag_debug_module_grant_vector)) OR (or_reduce(nios2_fast_fpu_jtag_debug_module_grant_vector))) OR (or_reduce(nios2_fast_fpu_jtag_debug_module_grant_vector))) OR (or_reduce(nios2_fast_fpu_jtag_debug_module_grant_vector));
  --nios2_fast_fpu_jtag_debug_module_end_xfer assignment, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_end_xfer <= NOT ((nios2_fast_fpu_jtag_debug_module_waits_for_read OR nios2_fast_fpu_jtag_debug_module_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_fast_fpu_jtag_debug_module arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_fast_fpu_jtag_debug_module <= nios2_fast_fpu_jtag_debug_module_end_xfer AND (((NOT nios2_fast_fpu_jtag_debug_module_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_fast_fpu_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_fast_fpu_jtag_debug_module AND nios2_fast_fpu_jtag_debug_module_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_fast_fpu_jtag_debug_module AND NOT nios2_fast_fpu_jtag_debug_module_non_bursting_master_requests));
  --nios2_fast_fpu_jtag_debug_module_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fast_fpu_jtag_debug_module_arb_share_counter <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fast_fpu_jtag_debug_module_arb_counter_enable) = '1' then 
        nios2_fast_fpu_jtag_debug_module_arb_share_counter <= nios2_fast_fpu_jtag_debug_module_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_fast_fpu_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fast_fpu_jtag_debug_module_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(nios2_fast_fpu_jtag_debug_module_master_qreq_vector) AND end_xfer_arb_share_counter_term_nios2_fast_fpu_jtag_debug_module)) OR ((end_xfer_arb_share_counter_term_nios2_fast_fpu_jtag_debug_module AND NOT nios2_fast_fpu_jtag_debug_module_non_bursting_master_requests)))) = '1' then 
        nios2_fast_fpu_jtag_debug_module_slavearbiterlockenable <= or_reduce(nios2_fast_fpu_jtag_debug_module_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --nios2_fpu_burst_4/downstream nios2_fast_fpu/jtag_debug_module arbiterlock, which is an e_assign
  nios2_fpu_burst_4_downstream_arbiterlock <= nios2_fast_fpu_jtag_debug_module_slavearbiterlockenable AND nios2_fpu_burst_4_downstream_continuerequest;
  --nios2_fast_fpu_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_slavearbiterlockenable2 <= or_reduce(nios2_fast_fpu_jtag_debug_module_arb_share_counter_next_value);
  --nios2_fpu_burst_4/downstream nios2_fast_fpu/jtag_debug_module arbiterlock2, which is an e_assign
  nios2_fpu_burst_4_downstream_arbiterlock2 <= nios2_fast_fpu_jtag_debug_module_slavearbiterlockenable2 AND nios2_fpu_burst_4_downstream_continuerequest;
  --nios2_fpu_burst_5/downstream nios2_fast_fpu/jtag_debug_module arbiterlock, which is an e_assign
  nios2_fpu_burst_5_downstream_arbiterlock <= nios2_fast_fpu_jtag_debug_module_slavearbiterlockenable AND nios2_fpu_burst_5_downstream_continuerequest;
  --nios2_fpu_burst_5/downstream nios2_fast_fpu/jtag_debug_module arbiterlock2, which is an e_assign
  nios2_fpu_burst_5_downstream_arbiterlock2 <= nios2_fast_fpu_jtag_debug_module_slavearbiterlockenable2 AND nios2_fpu_burst_5_downstream_continuerequest;
  --nios2_fpu_burst_5/downstream granted nios2_fast_fpu/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_nios2_fpu_burst_5_downstream_granted_slave_nios2_fast_fpu_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_nios2_fpu_burst_5_downstream_granted_slave_nios2_fast_fpu_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_5_downstream_saved_grant_nios2_fast_fpu_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_jtag_debug_module_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_5_downstream_granted_slave_nios2_fast_fpu_jtag_debug_module))))));
    end if;

  end process;

  --nios2_fpu_burst_5_downstream_continuerequest continued request, which is an e_mux
  nios2_fpu_burst_5_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_5_downstream_granted_slave_nios2_fast_fpu_jtag_debug_module))) AND std_logic_vector'("00000000000000000000000000000001")));
  --nios2_fast_fpu_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  nios2_fast_fpu_jtag_debug_module_any_continuerequest <= nios2_fpu_burst_5_downstream_continuerequest OR nios2_fpu_burst_4_downstream_continuerequest;
  internal_nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module <= internal_nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module AND NOT ((((nios2_fpu_burst_4_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_4_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000")))))) OR nios2_fpu_burst_5_downstream_arbiterlock));
  --local readdatavalid nios2_fpu_burst_4_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module, which is an e_mux
  nios2_fpu_burst_4_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module <= (internal_nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module AND nios2_fpu_burst_4_downstream_read) AND NOT nios2_fast_fpu_jtag_debug_module_waits_for_read;
  --nios2_fast_fpu_jtag_debug_module_writedata mux, which is an e_mux
  nios2_fast_fpu_jtag_debug_module_writedata <= A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module)) = '1'), nios2_fpu_burst_4_downstream_writedata, nios2_fpu_burst_5_downstream_writedata);
  internal_nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_5_downstream_read OR nios2_fpu_burst_5_downstream_write)))))));
  --nios2_fpu_burst_4/downstream granted nios2_fast_fpu/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_nios2_fpu_burst_4_downstream_granted_slave_nios2_fast_fpu_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_nios2_fpu_burst_4_downstream_granted_slave_nios2_fast_fpu_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_4_downstream_saved_grant_nios2_fast_fpu_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_jtag_debug_module_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_4_downstream_granted_slave_nios2_fast_fpu_jtag_debug_module))))));
    end if;

  end process;

  --nios2_fpu_burst_4_downstream_continuerequest continued request, which is an e_mux
  nios2_fpu_burst_4_downstream_continuerequest <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_4_downstream_granted_slave_nios2_fast_fpu_jtag_debug_module))) AND std_logic_vector'("00000000000000000000000000000001")));
  internal_nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module <= internal_nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module AND NOT ((((nios2_fpu_burst_5_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_5_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000")))))) OR nios2_fpu_burst_4_downstream_arbiterlock));
  --local readdatavalid nios2_fpu_burst_5_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module, which is an e_mux
  nios2_fpu_burst_5_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module <= (internal_nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module AND nios2_fpu_burst_5_downstream_read) AND NOT nios2_fast_fpu_jtag_debug_module_waits_for_read;
  --allow new arb cycle for nios2_fast_fpu/jtag_debug_module, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_allow_new_arb_cycle <= NOT nios2_fpu_burst_4_downstream_arbiterlock AND NOT nios2_fpu_burst_5_downstream_arbiterlock;
  --nios2_fpu_burst_5/downstream assignment into master qualified-requests vector for nios2_fast_fpu/jtag_debug_module, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_master_qreq_vector(0) <= internal_nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module;
  --nios2_fpu_burst_5/downstream grant nios2_fast_fpu/jtag_debug_module, which is an e_assign
  internal_nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module <= nios2_fast_fpu_jtag_debug_module_grant_vector(0);
  --nios2_fpu_burst_5/downstream saved-grant nios2_fast_fpu/jtag_debug_module, which is an e_assign
  nios2_fpu_burst_5_downstream_saved_grant_nios2_fast_fpu_jtag_debug_module <= nios2_fast_fpu_jtag_debug_module_arb_winner(0);
  --nios2_fpu_burst_4/downstream assignment into master qualified-requests vector for nios2_fast_fpu/jtag_debug_module, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_master_qreq_vector(1) <= internal_nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module;
  --nios2_fpu_burst_4/downstream grant nios2_fast_fpu/jtag_debug_module, which is an e_assign
  internal_nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module <= nios2_fast_fpu_jtag_debug_module_grant_vector(1);
  --nios2_fpu_burst_4/downstream saved-grant nios2_fast_fpu/jtag_debug_module, which is an e_assign
  nios2_fpu_burst_4_downstream_saved_grant_nios2_fast_fpu_jtag_debug_module <= nios2_fast_fpu_jtag_debug_module_arb_winner(1);
  --nios2_fast_fpu/jtag_debug_module chosen-master double-vector, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((nios2_fast_fpu_jtag_debug_module_master_qreq_vector & nios2_fast_fpu_jtag_debug_module_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT nios2_fast_fpu_jtag_debug_module_master_qreq_vector & NOT nios2_fast_fpu_jtag_debug_module_master_qreq_vector))) + (std_logic_vector'("000") & (nios2_fast_fpu_jtag_debug_module_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  nios2_fast_fpu_jtag_debug_module_arb_winner <= A_WE_StdLogicVector((std_logic'(((nios2_fast_fpu_jtag_debug_module_allow_new_arb_cycle AND or_reduce(nios2_fast_fpu_jtag_debug_module_grant_vector)))) = '1'), nios2_fast_fpu_jtag_debug_module_grant_vector, nios2_fast_fpu_jtag_debug_module_saved_chosen_master_vector);
  --saved nios2_fast_fpu_jtag_debug_module_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fast_fpu_jtag_debug_module_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fast_fpu_jtag_debug_module_allow_new_arb_cycle) = '1' then 
        nios2_fast_fpu_jtag_debug_module_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(nios2_fast_fpu_jtag_debug_module_grant_vector)) = '1'), nios2_fast_fpu_jtag_debug_module_grant_vector, nios2_fast_fpu_jtag_debug_module_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  nios2_fast_fpu_jtag_debug_module_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((nios2_fast_fpu_jtag_debug_module_chosen_master_double_vector(1) OR nios2_fast_fpu_jtag_debug_module_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((nios2_fast_fpu_jtag_debug_module_chosen_master_double_vector(0) OR nios2_fast_fpu_jtag_debug_module_chosen_master_double_vector(2)))));
  --nios2_fast_fpu/jtag_debug_module chosen master rotated left, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(nios2_fast_fpu_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(nios2_fast_fpu_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --nios2_fast_fpu/jtag_debug_module's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fast_fpu_jtag_debug_module_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(nios2_fast_fpu_jtag_debug_module_grant_vector)) = '1' then 
        nios2_fast_fpu_jtag_debug_module_arb_addend <= A_WE_StdLogicVector((std_logic'(nios2_fast_fpu_jtag_debug_module_end_xfer) = '1'), nios2_fast_fpu_jtag_debug_module_chosen_master_rot_left, nios2_fast_fpu_jtag_debug_module_grant_vector);
      end if;
    end if;

  end process;

  nios2_fast_fpu_jtag_debug_module_begintransfer <= nios2_fast_fpu_jtag_debug_module_begins_xfer;
  --assign nios2_fast_fpu_jtag_debug_module_resetrequest_from_sa = nios2_fast_fpu_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_resetrequest_from_sa <= nios2_fast_fpu_jtag_debug_module_resetrequest;
  nios2_fast_fpu_jtag_debug_module_chipselect <= internal_nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module OR internal_nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module;
  --nios2_fast_fpu_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_fast_fpu_jtag_debug_module_begins_xfer) = '1'), nios2_fast_fpu_jtag_debug_module_unreg_firsttransfer, nios2_fast_fpu_jtag_debug_module_reg_firsttransfer);
  --nios2_fast_fpu_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_unreg_firsttransfer <= NOT ((nios2_fast_fpu_jtag_debug_module_slavearbiterlockenable AND nios2_fast_fpu_jtag_debug_module_any_continuerequest));
  --nios2_fast_fpu_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fast_fpu_jtag_debug_module_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fast_fpu_jtag_debug_module_begins_xfer) = '1' then 
        nios2_fast_fpu_jtag_debug_module_reg_firsttransfer <= nios2_fast_fpu_jtag_debug_module_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_fast_fpu_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_beginbursttransfer_internal <= nios2_fast_fpu_jtag_debug_module_begins_xfer;
  --nios2_fast_fpu_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_arbitration_holdoff_internal <= nios2_fast_fpu_jtag_debug_module_begins_xfer AND nios2_fast_fpu_jtag_debug_module_firsttransfer;
  --nios2_fast_fpu_jtag_debug_module_write assignment, which is an e_mux
  nios2_fast_fpu_jtag_debug_module_write <= ((internal_nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module AND nios2_fpu_burst_4_downstream_write)) OR ((internal_nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module AND nios2_fpu_burst_5_downstream_write));
  shifted_address_to_nios2_fast_fpu_jtag_debug_module_from_nios2_fpu_burst_4_downstream <= nios2_fpu_burst_4_downstream_address_to_slave;
  --nios2_fast_fpu_jtag_debug_module_address mux, which is an e_mux
  nios2_fast_fpu_jtag_debug_module_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module)) = '1'), (A_SRL(shifted_address_to_nios2_fast_fpu_jtag_debug_module_from_nios2_fpu_burst_4_downstream,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_nios2_fast_fpu_jtag_debug_module_from_nios2_fpu_burst_5_downstream,std_logic_vector'("00000000000000000000000000000010")))), 9);
  shifted_address_to_nios2_fast_fpu_jtag_debug_module_from_nios2_fpu_burst_5_downstream <= nios2_fpu_burst_5_downstream_address_to_slave;
  --d1_nios2_fast_fpu_jtag_debug_module_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_fast_fpu_jtag_debug_module_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_fast_fpu_jtag_debug_module_end_xfer <= nios2_fast_fpu_jtag_debug_module_end_xfer;
    end if;

  end process;

  --nios2_fast_fpu_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  nios2_fast_fpu_jtag_debug_module_waits_for_read <= nios2_fast_fpu_jtag_debug_module_in_a_read_cycle AND nios2_fast_fpu_jtag_debug_module_begins_xfer;
  --nios2_fast_fpu_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_in_a_read_cycle <= ((internal_nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module AND nios2_fpu_burst_4_downstream_read)) OR ((internal_nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module AND nios2_fpu_burst_5_downstream_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_fast_fpu_jtag_debug_module_in_a_read_cycle;
  --nios2_fast_fpu_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  nios2_fast_fpu_jtag_debug_module_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_jtag_debug_module_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --nios2_fast_fpu_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  nios2_fast_fpu_jtag_debug_module_in_a_write_cycle <= ((internal_nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module AND nios2_fpu_burst_4_downstream_write)) OR ((internal_nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module AND nios2_fpu_burst_5_downstream_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_fast_fpu_jtag_debug_module_in_a_write_cycle;
  wait_for_nios2_fast_fpu_jtag_debug_module_counter <= std_logic'('0');
  --nios2_fast_fpu_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  nios2_fast_fpu_jtag_debug_module_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_4_downstream_byteenable)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_5_downstream_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))), 4);
  --debugaccess mux, which is an e_mux
  nios2_fast_fpu_jtag_debug_module_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_4_downstream_debugaccess))), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_5_downstream_debugaccess))), std_logic_vector'("00000000000000000000000000000000"))));
  --vhdl renameroo for output signals
  nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module <= internal_nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module;
  --vhdl renameroo for output signals
  nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module <= internal_nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module;
  --vhdl renameroo for output signals
  nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module <= internal_nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module;
  --vhdl renameroo for output signals
  nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module <= internal_nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module;
  --vhdl renameroo for output signals
  nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module <= internal_nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module;
  --vhdl renameroo for output signals
  nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module <= internal_nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module;
--synthesis translate_off
    --nios2_fast_fpu/jtag_debug_module enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --nios2_fpu_burst_4/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line11 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_4_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line11, now);
          write(write_line11, string'(": "));
          write(write_line11, string'("nios2_fpu_burst_4/downstream drove 0 on its 'arbitrationshare' port while accessing slave nios2_fast_fpu/jtag_debug_module"));
          write(output, write_line11.all);
          deallocate (write_line11);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_4/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line12 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_4_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line12, now);
          write(write_line12, string'(": "));
          write(write_line12, string'("nios2_fpu_burst_4/downstream drove 0 on its 'burstcount' port while accessing slave nios2_fast_fpu/jtag_debug_module"));
          write(output, write_line12.all);
          deallocate (write_line12);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_5/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line13 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_5_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line13, now);
          write(write_line13, string'(": "));
          write(write_line13, string'("nios2_fpu_burst_5/downstream drove 0 on its 'arbitrationshare' port while accessing slave nios2_fast_fpu/jtag_debug_module"));
          write(output, write_line13.all);
          deallocate (write_line13);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_5/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line14 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_5_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line14, now);
          write(write_line14, string'(": "));
          write(write_line14, string'("nios2_fpu_burst_5/downstream drove 0 on its 'burstcount' port while accessing slave nios2_fast_fpu/jtag_debug_module"));
          write(output, write_line14.all);
          deallocate (write_line14);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line15 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line15, now);
          write(write_line15, string'(": "));
          write(write_line15, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line15.all);
          deallocate (write_line15);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line16 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_4_downstream_saved_grant_nios2_fast_fpu_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_5_downstream_saved_grant_nios2_fast_fpu_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line16, now);
          write(write_line16, string'(": "));
          write(write_line16, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line16.all);
          deallocate (write_line16);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_fast_fpu_custom_instruction_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fast_fpu_custom_instruction_master_multi_n : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_fast_fpu_custom_instruction_master_multi_start : IN STD_LOGIC;
                 signal nios2_fast_fpu_fpoint_s1_done_from_sa : IN STD_LOGIC;
                 signal nios2_fast_fpu_fpoint_s1_result_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done_from_sa : IN STD_LOGIC;
                 signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_fast_fpu_custom_instruction_master_multi_done : OUT STD_LOGIC;
                 signal nios2_fast_fpu_custom_instruction_master_multi_result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_custom_instruction_master_reset_n : OUT STD_LOGIC;
                 signal nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_fpoint_s1 : OUT STD_LOGIC;
                 signal nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0 : OUT STD_LOGIC;
                 signal nios2_fast_fpu_fpoint_s1_select : OUT STD_LOGIC;
                 signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select : OUT STD_LOGIC
              );
end entity nios2_fast_fpu_custom_instruction_master_arbitrator;


architecture europa of nios2_fast_fpu_custom_instruction_master_arbitrator is
                signal internal_nios2_fast_fpu_fpoint_s1_select :  STD_LOGIC;
                signal internal_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select :  STD_LOGIC;

begin

  internal_nios2_fast_fpu_fpoint_s1_select <= to_std_logic((Std_Logic_Vector'(nios2_fast_fpu_custom_instruction_master_multi_n(7 DOWNTO 2) & std_logic_vector'("00")) = std_logic_vector'("11111100")));
  internal_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select <= to_std_logic((Std_Logic_Vector'(nios2_fast_fpu_custom_instruction_master_multi_n(7 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("00000000")));
  nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_fpoint_s1 <= internal_nios2_fast_fpu_fpoint_s1_select AND nios2_fast_fpu_custom_instruction_master_multi_start;
  nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0 <= internal_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select AND nios2_fast_fpu_custom_instruction_master_multi_start;
  --nios2_fast_fpu_custom_instruction_master_multi_result mux, which is an e_mux
  nios2_fast_fpu_custom_instruction_master_multi_result <= ((A_REP(internal_nios2_fast_fpu_fpoint_s1_select, 32) AND nios2_fast_fpu_fpoint_s1_result_from_sa)) OR ((A_REP(internal_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select, 32) AND nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result_from_sa));
  --multi_done mux, which is an e_mux
  nios2_fast_fpu_custom_instruction_master_multi_done <= ((internal_nios2_fast_fpu_fpoint_s1_select AND nios2_fast_fpu_fpoint_s1_done_from_sa)) OR ((internal_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select AND nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done_from_sa));
  --nios2_fast_fpu_custom_instruction_master_reset_n local reset_n, which is an e_assign
  nios2_fast_fpu_custom_instruction_master_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_fast_fpu_fpoint_s1_select <= internal_nios2_fast_fpu_fpoint_s1_select;
  --vhdl renameroo for output signals
  nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select <= internal_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module;


architecture europa of jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity mmcdma_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity mmcdma_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module;


architecture europa of mmcdma_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity psw_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity psw_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module;


architecture europa of psw_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity spu_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity spu_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module;


architecture europa of spu_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity systimer_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity systimer_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module;


architecture europa of systimer_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sysuart_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity sysuart_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module;


architecture europa of sysuart_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity vga_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity vga_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module;


architecture europa of vga_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fast_fpu_data_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal core_clk : IN STD_LOGIC;
                 signal core_clk_reset_n : IN STD_LOGIC;
                 signal d1_nios2_fpu_burst_2_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_fpu_burst_5_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_fpu_burst_6_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_fpu_burst_8_upstream_end_xfer : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                 signal mmcdma_s1_irq_from_sa : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_address : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_write : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_2_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_2_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_fpu_burst_5_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_5_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_fpu_burst_6_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_6_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_fpu_burst_8_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_8_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal psw_s1_irq_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal spu_s1_irq_from_sa : IN STD_LOGIC;
                 signal systimer_s1_irq_from_sa : IN STD_LOGIC;
                 signal sysuart_s1_irq_from_sa : IN STD_LOGIC;
                 signal vga_s1_irq_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal nios2_fast_fpu_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_latency_counter : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_readdatavalid : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_waitrequest : OUT STD_LOGIC
              );
end entity nios2_fast_fpu_data_master_arbitrator;


architecture europa of nios2_fast_fpu_data_master_arbitrator is
component jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module;

component mmcdma_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component mmcdma_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module;

component psw_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component psw_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module;

component spu_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component spu_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module;

component systimer_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component systimer_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module;

component sysuart_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component sysuart_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module;

component vga_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component vga_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module;

                signal active_and_waiting_last_time :  STD_LOGIC;
                signal core_clk_jtag_uart_avalon_jtag_slave_irq_from_sa :  STD_LOGIC;
                signal core_clk_mmcdma_s1_irq_from_sa :  STD_LOGIC;
                signal core_clk_psw_s1_irq_from_sa :  STD_LOGIC;
                signal core_clk_spu_s1_irq_from_sa :  STD_LOGIC;
                signal core_clk_systimer_s1_irq_from_sa :  STD_LOGIC;
                signal core_clk_sysuart_s1_irq_from_sa :  STD_LOGIC;
                signal core_clk_vga_s1_irq_from_sa :  STD_LOGIC;
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dbs_rdv_count_enable :  STD_LOGIC;
                signal dbs_rdv_counter_overflow :  STD_LOGIC;
                signal internal_nios2_fast_fpu_data_master_address_to_slave :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal internal_nios2_fast_fpu_data_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_nios2_fast_fpu_data_master_latency_counter :  STD_LOGIC;
                signal internal_nios2_fast_fpu_data_master_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_data_master_address_last_time :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal nios2_fast_fpu_data_master_burstcount_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fast_fpu_data_master_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fast_fpu_data_master_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_data_master_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_data_master_dbs_rdv_counter_inc :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_data_master_is_granted_some_slave :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_next_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_data_master_read_but_no_slave_selected :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_read_last_time :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_run :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_write_last_time :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_nios2_fast_fpu_data_master_latency_counter :  STD_LOGIC;
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal pre_flush_nios2_fast_fpu_data_master_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream OR NOT nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream OR NOT nios2_fast_fpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_2_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream OR NOT nios2_fast_fpu_data_master_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_2_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_nios2_fast_fpu_data_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream OR NOT nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream OR NOT ((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_5_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream OR NOT ((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_5_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream OR NOT nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream OR NOT ((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_6_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream OR NOT ((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_6_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream OR NOT nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream OR NOT ((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_8_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream OR NOT ((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_8_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_fast_fpu_data_master_run <= r_1;
  --jtag_uart_avalon_jtag_slave_irq_from_sa from peri_clk to core_clk
  jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master : jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module
    port map(
      data_out => core_clk_jtag_uart_avalon_jtag_slave_irq_from_sa,
      clk => core_clk,
      data_in => jtag_uart_avalon_jtag_slave_irq_from_sa,
      reset_n => core_clk_reset_n
    );


  --irq assign, which is an e_assign
  nios2_fast_fpu_data_master_irq <= Std_Logic_Vector'(A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(core_clk_psw_s1_irq_from_sa) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(core_clk_jtag_uart_avalon_jtag_slave_irq_from_sa) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(core_clk_sysuart_s1_irq_from_sa) & A_ToStdLogicVector(core_clk_spu_s1_irq_from_sa) & A_ToStdLogicVector(core_clk_mmcdma_s1_irq_from_sa) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(core_clk_vga_s1_irq_from_sa) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(core_clk_systimer_s1_irq_from_sa));
  --mmcdma_s1_irq_from_sa from peri_clk to core_clk
  mmcdma_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master : mmcdma_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module
    port map(
      data_out => core_clk_mmcdma_s1_irq_from_sa,
      clk => core_clk,
      data_in => mmcdma_s1_irq_from_sa,
      reset_n => core_clk_reset_n
    );


  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_fast_fpu_data_master_address_to_slave <= nios2_fast_fpu_data_master_address(28 DOWNTO 0);
  --nios2_fast_fpu_data_master_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fast_fpu_data_master_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      nios2_fast_fpu_data_master_read_but_no_slave_selected <= (nios2_fast_fpu_data_master_read AND nios2_fast_fpu_data_master_run) AND NOT nios2_fast_fpu_data_master_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  nios2_fast_fpu_data_master_is_granted_some_slave <= ((nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream OR nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream) OR nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream) OR nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_nios2_fast_fpu_data_master_readdatavalid <= ((((nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream AND dbs_rdv_counter_overflow)) OR nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream) OR nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream) OR nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream;
  --latent slave read data valid which is not flushed, which is an e_mux
  nios2_fast_fpu_data_master_readdatavalid <= ((((((nios2_fast_fpu_data_master_read_but_no_slave_selected OR pre_flush_nios2_fast_fpu_data_master_readdatavalid) OR nios2_fast_fpu_data_master_read_but_no_slave_selected) OR pre_flush_nios2_fast_fpu_data_master_readdatavalid) OR nios2_fast_fpu_data_master_read_but_no_slave_selected) OR pre_flush_nios2_fast_fpu_data_master_readdatavalid) OR nios2_fast_fpu_data_master_read_but_no_slave_selected) OR pre_flush_nios2_fast_fpu_data_master_readdatavalid;
  --input to latent dbs-16 stored 0, which is an e_mux
  p1_dbs_latent_16_reg_segment_0 <= nios2_fpu_burst_2_upstream_readdata_from_sa;
  --dbs register for latent dbs-16 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_16_reg_segment_0 <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((nios2_fast_fpu_data_master_dbs_rdv_counter(1))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
      end if;
    end if;

  end process;

  --nios2_fast_fpu/data_master readdata mux, which is an e_mux
  nios2_fast_fpu_data_master_readdata <= ((((A_REP(NOT nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream, 32) OR Std_Logic_Vector'(nios2_fpu_burst_2_upstream_readdata_from_sa(15 DOWNTO 0) & dbs_latent_16_reg_segment_0))) AND ((A_REP(NOT nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream, 32) OR nios2_fpu_burst_5_upstream_readdata_from_sa))) AND ((A_REP(NOT nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream, 32) OR nios2_fpu_burst_6_upstream_readdata_from_sa))) AND ((A_REP(NOT nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream, 32) OR nios2_fpu_burst_8_upstream_readdata_from_sa));
  --mux write dbs 1, which is an e_mux
  nios2_fast_fpu_data_master_dbs_write_16 <= A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_dbs_address(1))) = '1'), nios2_fast_fpu_data_master_writedata(31 DOWNTO 16), nios2_fast_fpu_data_master_writedata(15 DOWNTO 0));
  --actual waitrequest port, which is an e_assign
  internal_nios2_fast_fpu_data_master_waitrequest <= NOT nios2_fast_fpu_data_master_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_nios2_fast_fpu_data_master_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_nios2_fast_fpu_data_master_latency_counter <= p1_nios2_fast_fpu_data_master_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_nios2_fast_fpu_data_master_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((nios2_fast_fpu_data_master_run AND nios2_fast_fpu_data_master_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_nios2_fast_fpu_data_master_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --dbs count increment, which is an e_mux
  nios2_fast_fpu_data_master_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000000")), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_nios2_fast_fpu_data_master_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_nios2_fast_fpu_data_master_dbs_address)) + (std_logic_vector'("0") & (nios2_fast_fpu_data_master_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_nios2_fast_fpu_data_master_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_nios2_fast_fpu_data_master_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --p1 dbs rdv counter, which is an e_assign
  nios2_fast_fpu_data_master_next_dbs_rdv_counter <= A_EXT (((std_logic_vector'("0") & (nios2_fast_fpu_data_master_dbs_rdv_counter)) + (std_logic_vector'("0") & (nios2_fast_fpu_data_master_dbs_rdv_counter_inc))), 2);
  --nios2_fast_fpu_data_master_rdv_inc_mux, which is an e_mux
  nios2_fast_fpu_data_master_dbs_rdv_counter_inc <= std_logic_vector'("10");
  --master any slave rdv, which is an e_mux
  dbs_rdv_count_enable <= nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream;
  --dbs rdv counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fast_fpu_data_master_dbs_rdv_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_rdv_count_enable) = '1' then 
        nios2_fast_fpu_data_master_dbs_rdv_counter <= nios2_fast_fpu_data_master_next_dbs_rdv_counter;
      end if;
    end if;

  end process;

  --dbs rdv counter overflow, which is an e_assign
  dbs_rdv_counter_overflow <= nios2_fast_fpu_data_master_dbs_rdv_counter(1) AND NOT nios2_fast_fpu_data_master_next_dbs_rdv_counter(1);
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic(((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream AND nios2_fast_fpu_data_master_read)))) AND std_logic_vector'("00000000000000000000000000000000")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_2_upstream_waitrequest_from_sa))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream AND nios2_fast_fpu_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_2_upstream_waitrequest_from_sa)))))));
  --psw_s1_irq_from_sa from peri_clk to core_clk
  psw_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master : psw_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module
    port map(
      data_out => core_clk_psw_s1_irq_from_sa,
      clk => core_clk,
      data_in => psw_s1_irq_from_sa,
      reset_n => core_clk_reset_n
    );


  --spu_s1_irq_from_sa from peri_clk to core_clk
  spu_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master : spu_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module
    port map(
      data_out => core_clk_spu_s1_irq_from_sa,
      clk => core_clk,
      data_in => spu_s1_irq_from_sa,
      reset_n => core_clk_reset_n
    );


  --systimer_s1_irq_from_sa from peri_clk to core_clk
  systimer_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master : systimer_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module
    port map(
      data_out => core_clk_systimer_s1_irq_from_sa,
      clk => core_clk,
      data_in => systimer_s1_irq_from_sa,
      reset_n => core_clk_reset_n
    );


  --sysuart_s1_irq_from_sa from peri_clk to core_clk
  sysuart_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master : sysuart_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module
    port map(
      data_out => core_clk_sysuart_s1_irq_from_sa,
      clk => core_clk,
      data_in => sysuart_s1_irq_from_sa,
      reset_n => core_clk_reset_n
    );


  --vga_s1_irq_from_sa from peri_clk to core_clk
  vga_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master : vga_s1_irq_from_sa_clock_crossing_nios2_fast_fpu_data_master_module
    port map(
      data_out => core_clk_vga_s1_irq_from_sa,
      clk => core_clk,
      data_in => vga_s1_irq_from_sa,
      reset_n => core_clk_reset_n
    );


  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_address_to_slave <= internal_nios2_fast_fpu_data_master_address_to_slave;
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_dbs_address <= internal_nios2_fast_fpu_data_master_dbs_address;
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_latency_counter <= internal_nios2_fast_fpu_data_master_latency_counter;
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_waitrequest <= internal_nios2_fast_fpu_data_master_waitrequest;
--synthesis translate_off
    --nios2_fast_fpu_data_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fast_fpu_data_master_address_last_time <= std_logic_vector'("00000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fast_fpu_data_master_address_last_time <= nios2_fast_fpu_data_master_address;
      end if;

    end process;

    --nios2_fast_fpu/data_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_fast_fpu_data_master_waitrequest AND ((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write));
      end if;

    end process;

    --nios2_fast_fpu_data_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line17 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fast_fpu_data_master_address /= nios2_fast_fpu_data_master_address_last_time))))) = '1' then 
          write(write_line17, now);
          write(write_line17, string'(": "));
          write(write_line17, string'("nios2_fast_fpu_data_master_address did not heed wait!!!"));
          write(output, write_line17.all);
          deallocate (write_line17);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fast_fpu_data_master_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fast_fpu_data_master_burstcount_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_fast_fpu_data_master_burstcount_last_time <= nios2_fast_fpu_data_master_burstcount;
      end if;

    end process;

    --nios2_fast_fpu_data_master_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line18 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fast_fpu_data_master_burstcount /= nios2_fast_fpu_data_master_burstcount_last_time))))) = '1' then 
          write(write_line18, now);
          write(write_line18, string'(": "));
          write(write_line18, string'("nios2_fast_fpu_data_master_burstcount did not heed wait!!!"));
          write(output, write_line18.all);
          deallocate (write_line18);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fast_fpu_data_master_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fast_fpu_data_master_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_fast_fpu_data_master_byteenable_last_time <= nios2_fast_fpu_data_master_byteenable;
      end if;

    end process;

    --nios2_fast_fpu_data_master_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line19 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fast_fpu_data_master_byteenable /= nios2_fast_fpu_data_master_byteenable_last_time))))) = '1' then 
          write(write_line19, now);
          write(write_line19, string'(": "));
          write(write_line19, string'("nios2_fast_fpu_data_master_byteenable did not heed wait!!!"));
          write(output, write_line19.all);
          deallocate (write_line19);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fast_fpu_data_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fast_fpu_data_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fast_fpu_data_master_read_last_time <= nios2_fast_fpu_data_master_read;
      end if;

    end process;

    --nios2_fast_fpu_data_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line20 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fast_fpu_data_master_read) /= std_logic'(nios2_fast_fpu_data_master_read_last_time)))))) = '1' then 
          write(write_line20, now);
          write(write_line20, string'(": "));
          write(write_line20, string'("nios2_fast_fpu_data_master_read did not heed wait!!!"));
          write(output, write_line20.all);
          deallocate (write_line20);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fast_fpu_data_master_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fast_fpu_data_master_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fast_fpu_data_master_write_last_time <= nios2_fast_fpu_data_master_write;
      end if;

    end process;

    --nios2_fast_fpu_data_master_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line21 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fast_fpu_data_master_write) /= std_logic'(nios2_fast_fpu_data_master_write_last_time)))))) = '1' then 
          write(write_line21, now);
          write(write_line21, string'(": "));
          write(write_line21, string'("nios2_fast_fpu_data_master_write did not heed wait!!!"));
          write(output, write_line21.all);
          deallocate (write_line21);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fast_fpu_data_master_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fast_fpu_data_master_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fast_fpu_data_master_writedata_last_time <= nios2_fast_fpu_data_master_writedata;
      end if;

    end process;

    --nios2_fast_fpu_data_master_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line22 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_fast_fpu_data_master_writedata /= nios2_fast_fpu_data_master_writedata_last_time)))) AND nios2_fast_fpu_data_master_write)) = '1' then 
          write(write_line22, now);
          write(write_line22, string'(": "));
          write(write_line22, string'("nios2_fast_fpu_data_master_writedata did not heed wait!!!"));
          write(output, write_line22.all);
          deallocate (write_line22);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fast_fpu_instruction_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_nios2_fpu_burst_1_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_fpu_burst_4_upstream_end_xfer : IN STD_LOGIC;
                 signal d1_nios2_fpu_burst_7_upstream_end_xfer : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_address : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal nios2_fast_fpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_1_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_4_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal nios2_fpu_burst_7_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_7_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_fast_fpu_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal nios2_fast_fpu_instruction_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fast_fpu_instruction_master_latency_counter : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_instruction_master_readdatavalid : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_waitrequest : OUT STD_LOGIC
              );
end entity nios2_fast_fpu_instruction_master_arbitrator;


architecture europa of nios2_fast_fpu_instruction_master_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dbs_rdv_count_enable :  STD_LOGIC;
                signal dbs_rdv_counter_overflow :  STD_LOGIC;
                signal internal_nios2_fast_fpu_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal internal_nios2_fast_fpu_instruction_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_nios2_fast_fpu_instruction_master_latency_counter :  STD_LOGIC;
                signal internal_nios2_fast_fpu_instruction_master_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_instruction_master_address_last_time :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal nios2_fast_fpu_instruction_master_burstcount_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fast_fpu_instruction_master_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_instruction_master_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_instruction_master_dbs_rdv_counter_inc :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_instruction_master_is_granted_some_slave :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_next_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_instruction_master_read_but_no_slave_selected :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_read_last_time :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_run :  STD_LOGIC;
                signal p1_dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_nios2_fast_fpu_instruction_master_latency_counter :  STD_LOGIC;
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal pre_flush_nios2_fast_fpu_instruction_master_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream OR NOT nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream OR NOT nios2_fast_fpu_instruction_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_1_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_instruction_master_read)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream OR NOT nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream OR NOT (nios2_fast_fpu_instruction_master_read))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_4_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((nios2_fast_fpu_instruction_master_read))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream OR NOT nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream OR NOT (nios2_fast_fpu_instruction_master_read))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_7_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((nios2_fast_fpu_instruction_master_read))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_fast_fpu_instruction_master_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_fast_fpu_instruction_master_address_to_slave <= nios2_fast_fpu_instruction_master_address(27 DOWNTO 0);
  --nios2_fast_fpu_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fast_fpu_instruction_master_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      nios2_fast_fpu_instruction_master_read_but_no_slave_selected <= (nios2_fast_fpu_instruction_master_read AND nios2_fast_fpu_instruction_master_run) AND NOT nios2_fast_fpu_instruction_master_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  nios2_fast_fpu_instruction_master_is_granted_some_slave <= (nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream OR nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream) OR nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_nios2_fast_fpu_instruction_master_readdatavalid <= (((nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream AND dbs_rdv_counter_overflow)) OR nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream) OR nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream;
  --latent slave read data valid which is not flushed, which is an e_mux
  nios2_fast_fpu_instruction_master_readdatavalid <= ((((nios2_fast_fpu_instruction_master_read_but_no_slave_selected OR pre_flush_nios2_fast_fpu_instruction_master_readdatavalid) OR nios2_fast_fpu_instruction_master_read_but_no_slave_selected) OR pre_flush_nios2_fast_fpu_instruction_master_readdatavalid) OR nios2_fast_fpu_instruction_master_read_but_no_slave_selected) OR pre_flush_nios2_fast_fpu_instruction_master_readdatavalid;
  --input to latent dbs-16 stored 0, which is an e_mux
  p1_dbs_latent_16_reg_segment_0 <= nios2_fpu_burst_1_upstream_readdata_from_sa;
  --dbs register for latent dbs-16 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_16_reg_segment_0 <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((nios2_fast_fpu_instruction_master_dbs_rdv_counter(1))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
      end if;
    end if;

  end process;

  --nios2_fast_fpu/instruction_master readdata mux, which is an e_mux
  nios2_fast_fpu_instruction_master_readdata <= (((A_REP(NOT nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream, 32) OR Std_Logic_Vector'(nios2_fpu_burst_1_upstream_readdata_from_sa(15 DOWNTO 0) & dbs_latent_16_reg_segment_0))) AND ((A_REP(NOT nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream, 32) OR nios2_fpu_burst_4_upstream_readdata_from_sa))) AND ((A_REP(NOT nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream, 32) OR nios2_fpu_burst_7_upstream_readdata_from_sa));
  --actual waitrequest port, which is an e_assign
  internal_nios2_fast_fpu_instruction_master_waitrequest <= NOT nios2_fast_fpu_instruction_master_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_nios2_fast_fpu_instruction_master_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_nios2_fast_fpu_instruction_master_latency_counter <= p1_nios2_fast_fpu_instruction_master_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_nios2_fast_fpu_instruction_master_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((nios2_fast_fpu_instruction_master_run AND nios2_fast_fpu_instruction_master_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_instruction_master_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_nios2_fast_fpu_instruction_master_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --dbs count increment, which is an e_mux
  nios2_fast_fpu_instruction_master_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000000")), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_nios2_fast_fpu_instruction_master_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_nios2_fast_fpu_instruction_master_dbs_address)) + (std_logic_vector'("0") & (nios2_fast_fpu_instruction_master_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_nios2_fast_fpu_instruction_master_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_nios2_fast_fpu_instruction_master_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --p1 dbs rdv counter, which is an e_assign
  nios2_fast_fpu_instruction_master_next_dbs_rdv_counter <= A_EXT (((std_logic_vector'("0") & (nios2_fast_fpu_instruction_master_dbs_rdv_counter)) + (std_logic_vector'("0") & (nios2_fast_fpu_instruction_master_dbs_rdv_counter_inc))), 2);
  --nios2_fast_fpu_instruction_master_rdv_inc_mux, which is an e_mux
  nios2_fast_fpu_instruction_master_dbs_rdv_counter_inc <= std_logic_vector'("10");
  --master any slave rdv, which is an e_mux
  dbs_rdv_count_enable <= nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream;
  --dbs rdv counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fast_fpu_instruction_master_dbs_rdv_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_rdv_count_enable) = '1' then 
        nios2_fast_fpu_instruction_master_dbs_rdv_counter <= nios2_fast_fpu_instruction_master_next_dbs_rdv_counter;
      end if;
    end if;

  end process;

  --dbs rdv counter overflow, which is an e_assign
  dbs_rdv_counter_overflow <= nios2_fast_fpu_instruction_master_dbs_rdv_counter(1) AND NOT nios2_fast_fpu_instruction_master_next_dbs_rdv_counter(1);
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream AND nios2_fast_fpu_instruction_master_read)))) AND std_logic_vector'("00000000000000000000000000000000")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_1_upstream_waitrequest_from_sa)))));
  --vhdl renameroo for output signals
  nios2_fast_fpu_instruction_master_address_to_slave <= internal_nios2_fast_fpu_instruction_master_address_to_slave;
  --vhdl renameroo for output signals
  nios2_fast_fpu_instruction_master_dbs_address <= internal_nios2_fast_fpu_instruction_master_dbs_address;
  --vhdl renameroo for output signals
  nios2_fast_fpu_instruction_master_latency_counter <= internal_nios2_fast_fpu_instruction_master_latency_counter;
  --vhdl renameroo for output signals
  nios2_fast_fpu_instruction_master_waitrequest <= internal_nios2_fast_fpu_instruction_master_waitrequest;
--synthesis translate_off
    --nios2_fast_fpu_instruction_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fast_fpu_instruction_master_address_last_time <= std_logic_vector'("0000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fast_fpu_instruction_master_address_last_time <= nios2_fast_fpu_instruction_master_address;
      end if;

    end process;

    --nios2_fast_fpu/instruction_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_fast_fpu_instruction_master_waitrequest AND (nios2_fast_fpu_instruction_master_read);
      end if;

    end process;

    --nios2_fast_fpu_instruction_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line23 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fast_fpu_instruction_master_address /= nios2_fast_fpu_instruction_master_address_last_time))))) = '1' then 
          write(write_line23, now);
          write(write_line23, string'(": "));
          write(write_line23, string'("nios2_fast_fpu_instruction_master_address did not heed wait!!!"));
          write(output, write_line23.all);
          deallocate (write_line23);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fast_fpu_instruction_master_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fast_fpu_instruction_master_burstcount_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_fast_fpu_instruction_master_burstcount_last_time <= nios2_fast_fpu_instruction_master_burstcount;
      end if;

    end process;

    --nios2_fast_fpu_instruction_master_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line24 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fast_fpu_instruction_master_burstcount /= nios2_fast_fpu_instruction_master_burstcount_last_time))))) = '1' then 
          write(write_line24, now);
          write(write_line24, string'(": "));
          write(write_line24, string'("nios2_fast_fpu_instruction_master_burstcount did not heed wait!!!"));
          write(output, write_line24.all);
          deallocate (write_line24);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fast_fpu_instruction_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fast_fpu_instruction_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fast_fpu_instruction_master_read_last_time <= nios2_fast_fpu_instruction_master_read;
      end if;

    end process;

    --nios2_fast_fpu_instruction_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line25 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fast_fpu_instruction_master_read) /= std_logic'(nios2_fast_fpu_instruction_master_read_last_time)))))) = '1' then 
          write(write_line25, now);
          write(write_line25, string'(": "));
          write(write_line25, string'("nios2_fast_fpu_instruction_master_read did not heed wait!!!"));
          write(output, write_line25.all);
          deallocate (write_line25);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_fast_fpu_fpoint_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fast_fpu_custom_instruction_master_multi_clk_en : IN STD_LOGIC;
                 signal nios2_fast_fpu_custom_instruction_master_multi_dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_custom_instruction_master_multi_datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_custom_instruction_master_multi_n : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_fpoint_s1 : IN STD_LOGIC;
                 signal nios2_fast_fpu_fpoint_s1_done : IN STD_LOGIC;
                 signal nios2_fast_fpu_fpoint_s1_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_fpoint_s1_select : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_fast_fpu_fpoint_s1_clk_en : OUT STD_LOGIC;
                 signal nios2_fast_fpu_fpoint_s1_dataa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_fpoint_s1_datab : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_fpoint_s1_done_from_sa : OUT STD_LOGIC;
                 signal nios2_fast_fpu_fpoint_s1_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fast_fpu_fpoint_s1_reset : OUT STD_LOGIC;
                 signal nios2_fast_fpu_fpoint_s1_result_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_fpoint_s1_start : OUT STD_LOGIC
              );
end entity nios2_fast_fpu_fpoint_s1_arbitrator;


architecture europa of nios2_fast_fpu_fpoint_s1_arbitrator is

begin

  nios2_fast_fpu_fpoint_s1_clk_en <= nios2_fast_fpu_custom_instruction_master_multi_clk_en;
  nios2_fast_fpu_fpoint_s1_dataa <= nios2_fast_fpu_custom_instruction_master_multi_dataa;
  nios2_fast_fpu_fpoint_s1_datab <= nios2_fast_fpu_custom_instruction_master_multi_datab;
  nios2_fast_fpu_fpoint_s1_n <= nios2_fast_fpu_custom_instruction_master_multi_n (1 DOWNTO 0);
  nios2_fast_fpu_fpoint_s1_start <= nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_fpoint_s1;
  --assign nios2_fast_fpu_fpoint_s1_result_from_sa = nios2_fast_fpu_fpoint_s1_result so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fast_fpu_fpoint_s1_result_from_sa <= nios2_fast_fpu_fpoint_s1_result;
  --assign nios2_fast_fpu_fpoint_s1_done_from_sa = nios2_fast_fpu_fpoint_s1_done so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fast_fpu_fpoint_s1_done_from_sa <= nios2_fast_fpu_fpoint_s1_done;
  --nios2_fast_fpu_fpoint/s1 local reset_n, which is an e_assign
  nios2_fast_fpu_fpoint_s1_reset <= NOT reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fast_fpu_custom_instruction_master_multi_clk_en : IN STD_LOGIC;
                 signal nios2_fast_fpu_custom_instruction_master_multi_dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_custom_instruction_master_multi_datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_custom_instruction_master_multi_n : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0 : IN STD_LOGIC;
                 signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done : IN STD_LOGIC;
                 signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_clk_en : OUT STD_LOGIC;
                 signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_dataa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_datab : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done_from_sa : OUT STD_LOGIC;
                 signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_n : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_reset : OUT STD_LOGIC;
                 signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_start : OUT STD_LOGIC
              );
end entity nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_arbitrator;


architecture europa of nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_arbitrator is

begin

  nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_clk_en <= nios2_fast_fpu_custom_instruction_master_multi_clk_en;
  nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_dataa <= nios2_fast_fpu_custom_instruction_master_multi_dataa;
  nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_datab <= nios2_fast_fpu_custom_instruction_master_multi_datab;
  nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_n <= nios2_fast_fpu_custom_instruction_master_multi_n (2 DOWNTO 0);
  nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_start <= nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0;
  --assign nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result_from_sa = nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result_from_sa <= nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result;
  --assign nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done_from_sa = nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done_from_sa <= nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done;
  --nios2_fast_fpu_pixelsimd_inst/nios_custom_instruction_slave_0 local reset_n, which is an e_assign
  nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_reset <= NOT reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_nios2_fpu_burst_0_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_nios2_fpu_burst_0_upstream_module;


architecture europa of burstcount_fifo_for_nios2_fpu_burst_0_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_3 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_4 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_5 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_6 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_7 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal stage_8 :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_8;
  empty <= NOT(full_0);
  full_9 <= std_logic'('0');
  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic_vector'("00000000000");
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic_vector'("00000000000");
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic_vector'("00000000000");
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic_vector'("00000000000");
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic_vector'("00000000000");
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic_vector'("00000000000");
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("00000000000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("00000000000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("00000000000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 5);
  one_count_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 5);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_vga_m1_to_nios2_fpu_burst_0_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_vga_m1_to_nios2_fpu_burst_0_upstream_module;


architecture europa of rdv_fifo_for_vga_m1_to_nios2_fpu_burst_0_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_8;
  empty <= NOT(full_0);
  full_9 <= std_logic'('0');
  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 5);
  one_count_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 5);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_0_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_0_upstream_readdatavalid : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal vga_m1_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal vga_m1_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal vga_m1_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal vga_m1_latency_counter : IN STD_LOGIC;
                 signal vga_m1_read : IN STD_LOGIC;

              -- outputs:
                 signal d1_nios2_fpu_burst_0_upstream_end_xfer : OUT STD_LOGIC;
                 signal nios2_fpu_burst_0_upstream_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_0_upstream_burstcount : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal nios2_fpu_burst_0_upstream_byteaddress : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal nios2_fpu_burst_0_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fpu_burst_0_upstream_debugaccess : OUT STD_LOGIC;
                 signal nios2_fpu_burst_0_upstream_read : OUT STD_LOGIC;
                 signal nios2_fpu_burst_0_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_0_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_fpu_burst_0_upstream_write : OUT STD_LOGIC;
                 signal vga_m1_granted_nios2_fpu_burst_0_upstream : OUT STD_LOGIC;
                 signal vga_m1_qualified_request_nios2_fpu_burst_0_upstream : OUT STD_LOGIC;
                 signal vga_m1_read_data_valid_nios2_fpu_burst_0_upstream : OUT STD_LOGIC;
                 signal vga_m1_read_data_valid_nios2_fpu_burst_0_upstream_shift_register : OUT STD_LOGIC;
                 signal vga_m1_requests_nios2_fpu_burst_0_upstream : OUT STD_LOGIC
              );
end entity nios2_fpu_burst_0_upstream_arbitrator;


architecture europa of nios2_fpu_burst_0_upstream_arbitrator is
component burstcount_fifo_for_nios2_fpu_burst_0_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_nios2_fpu_burst_0_upstream_module;

component rdv_fifo_for_vga_m1_to_nios2_fpu_burst_0_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_vga_m1_to_nios2_fpu_burst_0_upstream_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_fpu_burst_0_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_fpu_burst_0_upstream_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal internal_nios2_fpu_burst_0_upstream_read :  STD_LOGIC;
                signal internal_nios2_fpu_burst_0_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_nios2_fpu_burst_0_upstream_write :  STD_LOGIC;
                signal internal_vga_m1_granted_nios2_fpu_burst_0_upstream :  STD_LOGIC;
                signal internal_vga_m1_qualified_request_nios2_fpu_burst_0_upstream :  STD_LOGIC;
                signal internal_vga_m1_requests_nios2_fpu_burst_0_upstream :  STD_LOGIC;
                signal module_input :  STD_LOGIC;
                signal module_input1 :  STD_LOGIC;
                signal module_input2 :  STD_LOGIC;
                signal module_input3 :  STD_LOGIC;
                signal module_input4 :  STD_LOGIC;
                signal module_input5 :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_allgrants :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_any_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_arb_counter_enable :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_arb_share_counter :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_begins_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_current_burst :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_end_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_grant_vector :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_in_a_read_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_in_a_write_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_load_fifo :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_master_qreq_vector :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_next_burst_count :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_reg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_selected_burstcount :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_waits_for_read :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_waits_for_write :  STD_LOGIC;
                signal p0_nios2_fpu_burst_0_upstream_load_fifo :  STD_LOGIC;
                signal vga_m1_arbiterlock :  STD_LOGIC;
                signal vga_m1_arbiterlock2 :  STD_LOGIC;
                signal vga_m1_continuerequest :  STD_LOGIC;
                signal vga_m1_rdv_fifo_empty_nios2_fpu_burst_0_upstream :  STD_LOGIC;
                signal vga_m1_rdv_fifo_output_from_nios2_fpu_burst_0_upstream :  STD_LOGIC;
                signal vga_m1_saved_grant_nios2_fpu_burst_0_upstream :  STD_LOGIC;
                signal wait_for_nios2_fpu_burst_0_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_fpu_burst_0_upstream_end_xfer;
    end if;

  end process;

  nios2_fpu_burst_0_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_vga_m1_qualified_request_nios2_fpu_burst_0_upstream);
  --assign nios2_fpu_burst_0_upstream_readdata_from_sa = nios2_fpu_burst_0_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_0_upstream_readdata_from_sa <= nios2_fpu_burst_0_upstream_readdata;
  internal_vga_m1_requests_nios2_fpu_burst_0_upstream <= ((to_std_logic(((Std_Logic_Vector'(vga_m1_address_to_slave(31 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("00000000000000000000000000000000")))) AND (vga_m1_read))) AND vga_m1_read;
  --assign nios2_fpu_burst_0_upstream_waitrequest_from_sa = nios2_fpu_burst_0_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_fpu_burst_0_upstream_waitrequest_from_sa <= nios2_fpu_burst_0_upstream_waitrequest;
  --assign nios2_fpu_burst_0_upstream_readdatavalid_from_sa = nios2_fpu_burst_0_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_0_upstream_readdatavalid_from_sa <= nios2_fpu_burst_0_upstream_readdatavalid;
  --nios2_fpu_burst_0_upstream_arb_share_counter set values, which is an e_mux
  nios2_fpu_burst_0_upstream_arb_share_set_values <= std_logic_vector'("000000000001");
  --nios2_fpu_burst_0_upstream_non_bursting_master_requests mux, which is an e_mux
  nios2_fpu_burst_0_upstream_non_bursting_master_requests <= std_logic'('0');
  --nios2_fpu_burst_0_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_fpu_burst_0_upstream_any_bursting_master_saved_grant <= vga_m1_saved_grant_nios2_fpu_burst_0_upstream;
  --nios2_fpu_burst_0_upstream_arb_share_counter_next_value assignment, which is an e_assign
  nios2_fpu_burst_0_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_0_upstream_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000") & (nios2_fpu_burst_0_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_fpu_burst_0_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000") & (nios2_fpu_burst_0_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 12);
  --nios2_fpu_burst_0_upstream_allgrants all slave grants, which is an e_mux
  nios2_fpu_burst_0_upstream_allgrants <= nios2_fpu_burst_0_upstream_grant_vector;
  --nios2_fpu_burst_0_upstream_end_xfer assignment, which is an e_assign
  nios2_fpu_burst_0_upstream_end_xfer <= NOT ((nios2_fpu_burst_0_upstream_waits_for_read OR nios2_fpu_burst_0_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_fpu_burst_0_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_fpu_burst_0_upstream <= nios2_fpu_burst_0_upstream_end_xfer AND (((NOT nios2_fpu_burst_0_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_fpu_burst_0_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_fpu_burst_0_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_fpu_burst_0_upstream AND nios2_fpu_burst_0_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_0_upstream AND NOT nios2_fpu_burst_0_upstream_non_bursting_master_requests));
  --nios2_fpu_burst_0_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_0_upstream_arb_share_counter <= std_logic_vector'("000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_0_upstream_arb_counter_enable) = '1' then 
        nios2_fpu_burst_0_upstream_arb_share_counter <= nios2_fpu_burst_0_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_0_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_0_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_fpu_burst_0_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_fpu_burst_0_upstream)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_0_upstream AND NOT nios2_fpu_burst_0_upstream_non_bursting_master_requests)))) = '1' then 
        nios2_fpu_burst_0_upstream_slavearbiterlockenable <= or_reduce(nios2_fpu_burst_0_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --vga/m1 nios2_fpu_burst_0/upstream arbiterlock, which is an e_assign
  vga_m1_arbiterlock <= nios2_fpu_burst_0_upstream_slavearbiterlockenable AND vga_m1_continuerequest;
  --nios2_fpu_burst_0_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_fpu_burst_0_upstream_slavearbiterlockenable2 <= or_reduce(nios2_fpu_burst_0_upstream_arb_share_counter_next_value);
  --vga/m1 nios2_fpu_burst_0/upstream arbiterlock2, which is an e_assign
  vga_m1_arbiterlock2 <= nios2_fpu_burst_0_upstream_slavearbiterlockenable2 AND vga_m1_continuerequest;
  --nios2_fpu_burst_0_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_fpu_burst_0_upstream_any_continuerequest <= std_logic'('1');
  --vga_m1_continuerequest continued request, which is an e_assign
  vga_m1_continuerequest <= std_logic'('1');
  internal_vga_m1_qualified_request_nios2_fpu_burst_0_upstream <= internal_vga_m1_requests_nios2_fpu_burst_0_upstream AND NOT ((vga_m1_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(vga_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(vga_m1_latency_counter))))))))));
  --unique name for nios2_fpu_burst_0_upstream_move_on_to_next_transaction, which is an e_assign
  nios2_fpu_burst_0_upstream_move_on_to_next_transaction <= nios2_fpu_burst_0_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_0_upstream_load_fifo;
  --the currently selected burstcount for nios2_fpu_burst_0_upstream, which is an e_mux
  nios2_fpu_burst_0_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_vga_m1_granted_nios2_fpu_burst_0_upstream)) = '1'), (std_logic_vector'("0000000000000000000000") & (vga_m1_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 11);
  --burstcount_fifo_for_nios2_fpu_burst_0_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_nios2_fpu_burst_0_upstream : burstcount_fifo_for_nios2_fpu_burst_0_upstream_module
    port map(
      data_out => nios2_fpu_burst_0_upstream_transaction_burst_count,
      empty => nios2_fpu_burst_0_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input,
      clk => clk,
      data_in => nios2_fpu_burst_0_upstream_selected_burstcount,
      read => nios2_fpu_burst_0_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input1,
      write => module_input2
    );

  module_input <= std_logic'('0');
  module_input1 <= std_logic'('0');
  module_input2 <= ((in_a_read_cycle AND NOT nios2_fpu_burst_0_upstream_waits_for_read) AND nios2_fpu_burst_0_upstream_load_fifo) AND NOT ((nios2_fpu_burst_0_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_0_upstream_burstcount_fifo_empty));

  --nios2_fpu_burst_0_upstream current burst minus one, which is an e_assign
  nios2_fpu_burst_0_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000") & (nios2_fpu_burst_0_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 11);
  --what to load in current_burst, for nios2_fpu_burst_0_upstream, which is an e_mux
  nios2_fpu_burst_0_upstream_next_burst_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_0_upstream_waits_for_read)) AND NOT nios2_fpu_burst_0_upstream_load_fifo))) = '1'), (nios2_fpu_burst_0_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_0_upstream_waits_for_read) AND nios2_fpu_burst_0_upstream_this_cycle_is_the_last_burst) AND nios2_fpu_burst_0_upstream_burstcount_fifo_empty))) = '1'), (nios2_fpu_burst_0_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'((nios2_fpu_burst_0_upstream_this_cycle_is_the_last_burst)) = '1'), (nios2_fpu_burst_0_upstream_transaction_burst_count & A_ToStdLogicVector(std_logic'('0'))), (std_logic_vector'("0") & (nios2_fpu_burst_0_upstream_current_burst_minus_one))))), 11);
  --the current burst count for nios2_fpu_burst_0_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_0_upstream_current_burst <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((nios2_fpu_burst_0_upstream_readdatavalid_from_sa OR ((NOT nios2_fpu_burst_0_upstream_load_fifo AND ((in_a_read_cycle AND NOT nios2_fpu_burst_0_upstream_waits_for_read)))))) = '1' then 
        nios2_fpu_burst_0_upstream_current_burst <= nios2_fpu_burst_0_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_nios2_fpu_burst_0_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT nios2_fpu_burst_0_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_0_upstream_waits_for_read)) AND nios2_fpu_burst_0_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_0_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_0_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_0_upstream_waits_for_read)) AND NOT nios2_fpu_burst_0_upstream_load_fifo) OR nios2_fpu_burst_0_upstream_this_cycle_is_the_last_burst)) = '1' then 
        nios2_fpu_burst_0_upstream_load_fifo <= p0_nios2_fpu_burst_0_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for nios2_fpu_burst_0_upstream, which is an e_assign
  nios2_fpu_burst_0_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(nios2_fpu_burst_0_upstream_current_burst_minus_one)) AND nios2_fpu_burst_0_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_vga_m1_to_nios2_fpu_burst_0_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_vga_m1_to_nios2_fpu_burst_0_upstream : rdv_fifo_for_vga_m1_to_nios2_fpu_burst_0_upstream_module
    port map(
      data_out => vga_m1_rdv_fifo_output_from_nios2_fpu_burst_0_upstream,
      empty => open,
      fifo_contains_ones_n => vga_m1_rdv_fifo_empty_nios2_fpu_burst_0_upstream,
      full => open,
      clear_fifo => module_input3,
      clk => clk,
      data_in => internal_vga_m1_granted_nios2_fpu_burst_0_upstream,
      read => nios2_fpu_burst_0_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input4,
      write => module_input5
    );

  module_input3 <= std_logic'('0');
  module_input4 <= std_logic'('0');
  module_input5 <= in_a_read_cycle AND NOT nios2_fpu_burst_0_upstream_waits_for_read;

  vga_m1_read_data_valid_nios2_fpu_burst_0_upstream_shift_register <= NOT vga_m1_rdv_fifo_empty_nios2_fpu_burst_0_upstream;
  --local readdatavalid vga_m1_read_data_valid_nios2_fpu_burst_0_upstream, which is an e_mux
  vga_m1_read_data_valid_nios2_fpu_burst_0_upstream <= nios2_fpu_burst_0_upstream_readdatavalid_from_sa;
  --byteaddress mux for nios2_fpu_burst_0/upstream, which is an e_mux
  nios2_fpu_burst_0_upstream_byteaddress <= vga_m1_address_to_slave (25 DOWNTO 0);
  --master is always granted when requested
  internal_vga_m1_granted_nios2_fpu_burst_0_upstream <= internal_vga_m1_qualified_request_nios2_fpu_burst_0_upstream;
  --vga/m1 saved-grant nios2_fpu_burst_0/upstream, which is an e_assign
  vga_m1_saved_grant_nios2_fpu_burst_0_upstream <= internal_vga_m1_requests_nios2_fpu_burst_0_upstream;
  --allow new arb cycle for nios2_fpu_burst_0/upstream, which is an e_assign
  nios2_fpu_burst_0_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_fpu_burst_0_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_fpu_burst_0_upstream_master_qreq_vector <= std_logic'('1');
  --nios2_fpu_burst_0_upstream_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_0_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_fpu_burst_0_upstream_begins_xfer) = '1'), nios2_fpu_burst_0_upstream_unreg_firsttransfer, nios2_fpu_burst_0_upstream_reg_firsttransfer);
  --nios2_fpu_burst_0_upstream_unreg_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_0_upstream_unreg_firsttransfer <= NOT ((nios2_fpu_burst_0_upstream_slavearbiterlockenable AND nios2_fpu_burst_0_upstream_any_continuerequest));
  --nios2_fpu_burst_0_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_0_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_0_upstream_begins_xfer) = '1' then 
        nios2_fpu_burst_0_upstream_reg_firsttransfer <= nios2_fpu_burst_0_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_0_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  nios2_fpu_burst_0_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_nios2_fpu_burst_0_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000") & (nios2_fpu_burst_0_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000") & (internal_nios2_fpu_burst_0_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_nios2_fpu_burst_0_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000") & (nios2_fpu_burst_0_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000") & (nios2_fpu_burst_0_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 9);
  --nios2_fpu_burst_0_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_0_upstream_bbt_burstcounter <= std_logic_vector'("000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_0_upstream_begins_xfer) = '1' then 
        nios2_fpu_burst_0_upstream_bbt_burstcounter <= nios2_fpu_burst_0_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_0_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_fpu_burst_0_upstream_beginbursttransfer_internal <= nios2_fpu_burst_0_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000") & (nios2_fpu_burst_0_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --nios2_fpu_burst_0_upstream_read assignment, which is an e_mux
  internal_nios2_fpu_burst_0_upstream_read <= internal_vga_m1_granted_nios2_fpu_burst_0_upstream AND vga_m1_read;
  --nios2_fpu_burst_0_upstream_write assignment, which is an e_mux
  internal_nios2_fpu_burst_0_upstream_write <= std_logic'('0');
  --nios2_fpu_burst_0_upstream_address mux, which is an e_mux
  nios2_fpu_burst_0_upstream_address <= A_EXT (Std_Logic_Vector'(A_SRL(vga_m1_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(vga_m1_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 25);
  --d1_nios2_fpu_burst_0_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_fpu_burst_0_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_fpu_burst_0_upstream_end_xfer <= nios2_fpu_burst_0_upstream_end_xfer;
    end if;

  end process;

  --nios2_fpu_burst_0_upstream_waits_for_read in a cycle, which is an e_mux
  nios2_fpu_burst_0_upstream_waits_for_read <= nios2_fpu_burst_0_upstream_in_a_read_cycle AND internal_nios2_fpu_burst_0_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_0_upstream_in_a_read_cycle assignment, which is an e_assign
  nios2_fpu_burst_0_upstream_in_a_read_cycle <= internal_vga_m1_granted_nios2_fpu_burst_0_upstream AND vga_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_fpu_burst_0_upstream_in_a_read_cycle;
  --nios2_fpu_burst_0_upstream_waits_for_write in a cycle, which is an e_mux
  nios2_fpu_burst_0_upstream_waits_for_write <= nios2_fpu_burst_0_upstream_in_a_write_cycle AND internal_nios2_fpu_burst_0_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_0_upstream_in_a_write_cycle assignment, which is an e_assign
  nios2_fpu_burst_0_upstream_in_a_write_cycle <= std_logic'('0');
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_fpu_burst_0_upstream_in_a_write_cycle;
  wait_for_nios2_fpu_burst_0_upstream_counter <= std_logic'('0');
  --nios2_fpu_burst_0_upstream_byteenable byte enable port mux, which is an e_mux
  nios2_fpu_burst_0_upstream_byteenable <= A_EXT (-SIGNED(std_logic_vector'("00000000000000000000000000000001")), 2);
  --burstcount mux, which is an e_mux
  internal_nios2_fpu_burst_0_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_vga_m1_granted_nios2_fpu_burst_0_upstream)) = '1'), (std_logic_vector'("0000000000000000000000") & (vga_m1_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 10);
  --debugaccess mux, which is an e_mux
  nios2_fpu_burst_0_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_fpu_burst_0_upstream_burstcount <= internal_nios2_fpu_burst_0_upstream_burstcount;
  --vhdl renameroo for output signals
  nios2_fpu_burst_0_upstream_read <= internal_nios2_fpu_burst_0_upstream_read;
  --vhdl renameroo for output signals
  nios2_fpu_burst_0_upstream_waitrequest_from_sa <= internal_nios2_fpu_burst_0_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  nios2_fpu_burst_0_upstream_write <= internal_nios2_fpu_burst_0_upstream_write;
  --vhdl renameroo for output signals
  vga_m1_granted_nios2_fpu_burst_0_upstream <= internal_vga_m1_granted_nios2_fpu_burst_0_upstream;
  --vhdl renameroo for output signals
  vga_m1_qualified_request_nios2_fpu_burst_0_upstream <= internal_vga_m1_qualified_request_nios2_fpu_burst_0_upstream;
  --vhdl renameroo for output signals
  vga_m1_requests_nios2_fpu_burst_0_upstream <= internal_vga_m1_requests_nios2_fpu_burst_0_upstream;
--synthesis translate_off
    --nios2_fpu_burst_0/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --vga/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line26 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_vga_m1_requests_nios2_fpu_burst_0_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000") & (vga_m1_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line26, now);
          write(write_line26, string'(": "));
          write(write_line26, string'("vga/m1 drove 0 on its 'burstcount' port while accessing slave nios2_fpu_burst_0/upstream"));
          write(output, write_line26.all);
          deallocate (write_line26);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_0_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_0_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fpu_burst_0_downstream_granted_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_qualified_request_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_requests_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal nios2_fpu_burst_0_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_0_downstream_latency_counter : OUT STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_0_downstream_readdatavalid : OUT STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_reset_n : OUT STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_waitrequest : OUT STD_LOGIC
              );
end entity nios2_fpu_burst_0_downstream_arbitrator;


architecture europa of nios2_fpu_burst_0_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_fpu_burst_0_downstream_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal internal_nios2_fpu_burst_0_downstream_latency_counter :  STD_LOGIC;
                signal internal_nios2_fpu_burst_0_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_address_last_time :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_0_downstream_burstcount_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fpu_burst_0_downstream_is_granted_some_slave :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_read_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_run :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_write_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_nios2_fpu_burst_0_downstream_latency_counter :  STD_LOGIC;
                signal pre_flush_nios2_fpu_burst_0_downstream_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_0_downstream_qualified_request_sdram_s1 OR NOT nios2_fpu_burst_0_downstream_requests_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_0_downstream_granted_sdram_s1 OR NOT nios2_fpu_burst_0_downstream_qualified_request_sdram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_0_downstream_qualified_request_sdram_s1 OR NOT ((nios2_fpu_burst_0_downstream_read OR nios2_fpu_burst_0_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_0_downstream_read OR nios2_fpu_burst_0_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_0_downstream_qualified_request_sdram_s1 OR NOT ((nios2_fpu_burst_0_downstream_read OR nios2_fpu_burst_0_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_0_downstream_read OR nios2_fpu_burst_0_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_fpu_burst_0_downstream_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_fpu_burst_0_downstream_address_to_slave <= nios2_fpu_burst_0_downstream_address;
  --nios2_fpu_burst_0_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_0_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      nios2_fpu_burst_0_downstream_read_but_no_slave_selected <= (nios2_fpu_burst_0_downstream_read AND nios2_fpu_burst_0_downstream_run) AND NOT nios2_fpu_burst_0_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  nios2_fpu_burst_0_downstream_is_granted_some_slave <= nios2_fpu_burst_0_downstream_granted_sdram_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_nios2_fpu_burst_0_downstream_readdatavalid <= nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  nios2_fpu_burst_0_downstream_readdatavalid <= nios2_fpu_burst_0_downstream_read_but_no_slave_selected OR pre_flush_nios2_fpu_burst_0_downstream_readdatavalid;
  --nios2_fpu_burst_0/downstream readdata mux, which is an e_mux
  nios2_fpu_burst_0_downstream_readdata <= sdram_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_fpu_burst_0_downstream_waitrequest <= NOT nios2_fpu_burst_0_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_nios2_fpu_burst_0_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_nios2_fpu_burst_0_downstream_latency_counter <= p1_nios2_fpu_burst_0_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_nios2_fpu_burst_0_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((nios2_fpu_burst_0_downstream_run AND nios2_fpu_burst_0_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_0_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_0_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --nios2_fpu_burst_0_downstream_reset_n assignment, which is an e_assign
  nios2_fpu_burst_0_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_fpu_burst_0_downstream_address_to_slave <= internal_nios2_fpu_burst_0_downstream_address_to_slave;
  --vhdl renameroo for output signals
  nios2_fpu_burst_0_downstream_latency_counter <= internal_nios2_fpu_burst_0_downstream_latency_counter;
  --vhdl renameroo for output signals
  nios2_fpu_burst_0_downstream_waitrequest <= internal_nios2_fpu_burst_0_downstream_waitrequest;
--synthesis translate_off
    --nios2_fpu_burst_0_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_0_downstream_address_last_time <= std_logic_vector'("0000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_0_downstream_address_last_time <= nios2_fpu_burst_0_downstream_address;
      end if;

    end process;

    --nios2_fpu_burst_0/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_fpu_burst_0_downstream_waitrequest AND ((nios2_fpu_burst_0_downstream_read OR nios2_fpu_burst_0_downstream_write));
      end if;

    end process;

    --nios2_fpu_burst_0_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line27 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_0_downstream_address /= nios2_fpu_burst_0_downstream_address_last_time))))) = '1' then 
          write(write_line27, now);
          write(write_line27, string'(": "));
          write(write_line27, string'("nios2_fpu_burst_0_downstream_address did not heed wait!!!"));
          write(output, write_line27.all);
          deallocate (write_line27);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_0_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_0_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_0_downstream_burstcount_last_time <= nios2_fpu_burst_0_downstream_burstcount;
      end if;

    end process;

    --nios2_fpu_burst_0_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line28 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_0_downstream_burstcount) /= std_logic'(nios2_fpu_burst_0_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line28, now);
          write(write_line28, string'(": "));
          write(write_line28, string'("nios2_fpu_burst_0_downstream_burstcount did not heed wait!!!"));
          write(output, write_line28.all);
          deallocate (write_line28);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_0_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_0_downstream_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_0_downstream_byteenable_last_time <= nios2_fpu_burst_0_downstream_byteenable;
      end if;

    end process;

    --nios2_fpu_burst_0_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line29 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_0_downstream_byteenable /= nios2_fpu_burst_0_downstream_byteenable_last_time))))) = '1' then 
          write(write_line29, now);
          write(write_line29, string'(": "));
          write(write_line29, string'("nios2_fpu_burst_0_downstream_byteenable did not heed wait!!!"));
          write(output, write_line29.all);
          deallocate (write_line29);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_0_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_0_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_0_downstream_read_last_time <= nios2_fpu_burst_0_downstream_read;
      end if;

    end process;

    --nios2_fpu_burst_0_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line30 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_0_downstream_read) /= std_logic'(nios2_fpu_burst_0_downstream_read_last_time)))))) = '1' then 
          write(write_line30, now);
          write(write_line30, string'(": "));
          write(write_line30, string'("nios2_fpu_burst_0_downstream_read did not heed wait!!!"));
          write(output, write_line30.all);
          deallocate (write_line30);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_0_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_0_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_0_downstream_write_last_time <= nios2_fpu_burst_0_downstream_write;
      end if;

    end process;

    --nios2_fpu_burst_0_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line31 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_0_downstream_write) /= std_logic'(nios2_fpu_burst_0_downstream_write_last_time)))))) = '1' then 
          write(write_line31, now);
          write(write_line31, string'(": "));
          write(write_line31, string'("nios2_fpu_burst_0_downstream_write did not heed wait!!!"));
          write(output, write_line31.all);
          deallocate (write_line31);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_0_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_0_downstream_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_0_downstream_writedata_last_time <= nios2_fpu_burst_0_downstream_writedata;
      end if;

    end process;

    --nios2_fpu_burst_0_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line32 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_0_downstream_writedata /= nios2_fpu_burst_0_downstream_writedata_last_time)))) AND nios2_fpu_burst_0_downstream_write)) = '1' then 
          write(write_line32, now);
          write(write_line32, string'(": "));
          write(write_line32, string'("nios2_fpu_burst_0_downstream_writedata did not heed wait!!!"));
          write(output, write_line32.all);
          deallocate (write_line32);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_nios2_fpu_burst_1_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_nios2_fpu_burst_1_upstream_module;


architecture europa of burstcount_fifo_for_nios2_fpu_burst_1_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_3 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_4 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_5 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_6 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_7 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_8 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_8;
  empty <= NOT(full_0);
  full_9 <= std_logic'('0');
  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic_vector'("00000");
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic_vector'("00000");
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic_vector'("00000");
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic_vector'("00000");
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic_vector'("00000");
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic_vector'("00000");
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("00000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("00000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("00000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 5);
  one_count_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 5);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_1_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_1_upstream_module;


architecture europa of rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_1_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_8;
  empty <= NOT(full_0);
  full_9 <= std_logic'('0');
  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 5);
  one_count_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 5);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_1_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal nios2_fast_fpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fast_fpu_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fast_fpu_instruction_master_latency_counter : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_1_upstream_readdatavalid : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_nios2_fpu_burst_1_upstream_end_xfer : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream : OUT STD_LOGIC;
                 signal nios2_fpu_burst_1_upstream_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_1_upstream_byteaddress : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal nios2_fpu_burst_1_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fpu_burst_1_upstream_debugaccess : OUT STD_LOGIC;
                 signal nios2_fpu_burst_1_upstream_read : OUT STD_LOGIC;
                 signal nios2_fpu_burst_1_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_1_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_fpu_burst_1_upstream_write : OUT STD_LOGIC
              );
end entity nios2_fpu_burst_1_upstream_arbitrator;


architecture europa of nios2_fpu_burst_1_upstream_arbitrator is
component burstcount_fifo_for_nios2_fpu_burst_1_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_nios2_fpu_burst_1_upstream_module;

component rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_1_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_1_upstream_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_fpu_burst_1_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream :  STD_LOGIC;
                signal internal_nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream :  STD_LOGIC;
                signal internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream :  STD_LOGIC;
                signal internal_nios2_fpu_burst_1_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal module_input10 :  STD_LOGIC;
                signal module_input11 :  STD_LOGIC;
                signal module_input6 :  STD_LOGIC;
                signal module_input7 :  STD_LOGIC;
                signal module_input8 :  STD_LOGIC;
                signal module_input9 :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_continuerequest :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_rdv_fifo_empty_nios2_fpu_burst_1_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_rdv_fifo_output_from_nios2_fpu_burst_1_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_saved_grant_nios2_fpu_burst_1_upstream :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_allgrants :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_any_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_arb_counter_enable :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_arb_share_counter :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_1_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_1_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_1_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_begins_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_current_burst :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fpu_burst_1_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fpu_burst_1_upstream_end_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_grant_vector :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_in_a_read_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_in_a_write_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_load_fifo :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_master_qreq_vector :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_next_burst_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fpu_burst_1_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_reg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_selected_burstcount :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fpu_burst_1_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fpu_burst_1_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_waits_for_read :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_waits_for_write :  STD_LOGIC;
                signal p0_nios2_fpu_burst_1_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_nios2_fpu_burst_1_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_fpu_burst_1_upstream_end_xfer;
    end if;

  end process;

  nios2_fpu_burst_1_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream);
  --assign nios2_fpu_burst_1_upstream_readdata_from_sa = nios2_fpu_burst_1_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_1_upstream_readdata_from_sa <= nios2_fpu_burst_1_upstream_readdata;
  internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream <= ((to_std_logic(((Std_Logic_Vector'(nios2_fast_fpu_instruction_master_address_to_slave(27 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("0000000000000000000000000000")))) AND (nios2_fast_fpu_instruction_master_read))) AND nios2_fast_fpu_instruction_master_read;
  --assign nios2_fpu_burst_1_upstream_waitrequest_from_sa = nios2_fpu_burst_1_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_fpu_burst_1_upstream_waitrequest_from_sa <= nios2_fpu_burst_1_upstream_waitrequest;
  --assign nios2_fpu_burst_1_upstream_readdatavalid_from_sa = nios2_fpu_burst_1_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_1_upstream_readdatavalid_from_sa <= nios2_fpu_burst_1_upstream_readdatavalid;
  --nios2_fpu_burst_1_upstream_arb_share_counter set values, which is an e_mux
  nios2_fpu_burst_1_upstream_arb_share_set_values <= std_logic_vector'("000001");
  --nios2_fpu_burst_1_upstream_non_bursting_master_requests mux, which is an e_mux
  nios2_fpu_burst_1_upstream_non_bursting_master_requests <= std_logic'('0');
  --nios2_fpu_burst_1_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_fpu_burst_1_upstream_any_bursting_master_saved_grant <= nios2_fast_fpu_instruction_master_saved_grant_nios2_fpu_burst_1_upstream;
  --nios2_fpu_burst_1_upstream_arb_share_counter_next_value assignment, which is an e_assign
  nios2_fpu_burst_1_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_1_upstream_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_1_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_fpu_burst_1_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_1_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 6);
  --nios2_fpu_burst_1_upstream_allgrants all slave grants, which is an e_mux
  nios2_fpu_burst_1_upstream_allgrants <= nios2_fpu_burst_1_upstream_grant_vector;
  --nios2_fpu_burst_1_upstream_end_xfer assignment, which is an e_assign
  nios2_fpu_burst_1_upstream_end_xfer <= NOT ((nios2_fpu_burst_1_upstream_waits_for_read OR nios2_fpu_burst_1_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_fpu_burst_1_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_fpu_burst_1_upstream <= nios2_fpu_burst_1_upstream_end_xfer AND (((NOT nios2_fpu_burst_1_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_fpu_burst_1_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_fpu_burst_1_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_fpu_burst_1_upstream AND nios2_fpu_burst_1_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_1_upstream AND NOT nios2_fpu_burst_1_upstream_non_bursting_master_requests));
  --nios2_fpu_burst_1_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_1_upstream_arb_share_counter <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_1_upstream_arb_counter_enable) = '1' then 
        nios2_fpu_burst_1_upstream_arb_share_counter <= nios2_fpu_burst_1_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_1_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_1_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_fpu_burst_1_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_fpu_burst_1_upstream)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_1_upstream AND NOT nios2_fpu_burst_1_upstream_non_bursting_master_requests)))) = '1' then 
        nios2_fpu_burst_1_upstream_slavearbiterlockenable <= or_reduce(nios2_fpu_burst_1_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --nios2_fast_fpu/instruction_master nios2_fpu_burst_1/upstream arbiterlock, which is an e_assign
  nios2_fast_fpu_instruction_master_arbiterlock <= nios2_fpu_burst_1_upstream_slavearbiterlockenable AND nios2_fast_fpu_instruction_master_continuerequest;
  --nios2_fpu_burst_1_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_fpu_burst_1_upstream_slavearbiterlockenable2 <= or_reduce(nios2_fpu_burst_1_upstream_arb_share_counter_next_value);
  --nios2_fast_fpu/instruction_master nios2_fpu_burst_1/upstream arbiterlock2, which is an e_assign
  nios2_fast_fpu_instruction_master_arbiterlock2 <= nios2_fpu_burst_1_upstream_slavearbiterlockenable2 AND nios2_fast_fpu_instruction_master_continuerequest;
  --nios2_fpu_burst_1_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_fpu_burst_1_upstream_any_continuerequest <= std_logic'('1');
  --nios2_fast_fpu_instruction_master_continuerequest continued request, which is an e_assign
  nios2_fast_fpu_instruction_master_continuerequest <= std_logic'('1');
  internal_nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream <= internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream AND NOT ((nios2_fast_fpu_instruction_master_read AND (((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_instruction_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_instruction_master_latency_counter))))))) OR (nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register)) OR (nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register)))));
  --unique name for nios2_fpu_burst_1_upstream_move_on_to_next_transaction, which is an e_assign
  nios2_fpu_burst_1_upstream_move_on_to_next_transaction <= nios2_fpu_burst_1_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_1_upstream_load_fifo;
  --the currently selected burstcount for nios2_fpu_burst_1_upstream, which is an e_mux
  nios2_fpu_burst_1_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_instruction_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 5);
  --burstcount_fifo_for_nios2_fpu_burst_1_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_nios2_fpu_burst_1_upstream : burstcount_fifo_for_nios2_fpu_burst_1_upstream_module
    port map(
      data_out => nios2_fpu_burst_1_upstream_transaction_burst_count,
      empty => nios2_fpu_burst_1_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input6,
      clk => clk,
      data_in => nios2_fpu_burst_1_upstream_selected_burstcount,
      read => nios2_fpu_burst_1_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input7,
      write => module_input8
    );

  module_input6 <= std_logic'('0');
  module_input7 <= std_logic'('0');
  module_input8 <= ((in_a_read_cycle AND NOT nios2_fpu_burst_1_upstream_waits_for_read) AND nios2_fpu_burst_1_upstream_load_fifo) AND NOT ((nios2_fpu_burst_1_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_1_upstream_burstcount_fifo_empty));

  --nios2_fpu_burst_1_upstream current burst minus one, which is an e_assign
  nios2_fpu_burst_1_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_1_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --what to load in current_burst, for nios2_fpu_burst_1_upstream, which is an e_mux
  nios2_fpu_burst_1_upstream_next_burst_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_1_upstream_waits_for_read)) AND NOT nios2_fpu_burst_1_upstream_load_fifo))) = '1'), (nios2_fpu_burst_1_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_1_upstream_waits_for_read) AND nios2_fpu_burst_1_upstream_this_cycle_is_the_last_burst) AND nios2_fpu_burst_1_upstream_burstcount_fifo_empty))) = '1'), (nios2_fpu_burst_1_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'((nios2_fpu_burst_1_upstream_this_cycle_is_the_last_burst)) = '1'), (nios2_fpu_burst_1_upstream_transaction_burst_count & A_ToStdLogicVector(std_logic'('0'))), (std_logic_vector'("0") & (nios2_fpu_burst_1_upstream_current_burst_minus_one))))), 5);
  --the current burst count for nios2_fpu_burst_1_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_1_upstream_current_burst <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((nios2_fpu_burst_1_upstream_readdatavalid_from_sa OR ((NOT nios2_fpu_burst_1_upstream_load_fifo AND ((in_a_read_cycle AND NOT nios2_fpu_burst_1_upstream_waits_for_read)))))) = '1' then 
        nios2_fpu_burst_1_upstream_current_burst <= nios2_fpu_burst_1_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_nios2_fpu_burst_1_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT nios2_fpu_burst_1_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_1_upstream_waits_for_read)) AND nios2_fpu_burst_1_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_1_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_1_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_1_upstream_waits_for_read)) AND NOT nios2_fpu_burst_1_upstream_load_fifo) OR nios2_fpu_burst_1_upstream_this_cycle_is_the_last_burst)) = '1' then 
        nios2_fpu_burst_1_upstream_load_fifo <= p0_nios2_fpu_burst_1_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for nios2_fpu_burst_1_upstream, which is an e_assign
  nios2_fpu_burst_1_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(nios2_fpu_burst_1_upstream_current_burst_minus_one)) AND nios2_fpu_burst_1_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_1_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_1_upstream : rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_1_upstream_module
    port map(
      data_out => nios2_fast_fpu_instruction_master_rdv_fifo_output_from_nios2_fpu_burst_1_upstream,
      empty => open,
      fifo_contains_ones_n => nios2_fast_fpu_instruction_master_rdv_fifo_empty_nios2_fpu_burst_1_upstream,
      full => open,
      clear_fifo => module_input9,
      clk => clk,
      data_in => internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream,
      read => nios2_fpu_burst_1_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input10,
      write => module_input11
    );

  module_input9 <= std_logic'('0');
  module_input10 <= std_logic'('0');
  module_input11 <= in_a_read_cycle AND NOT nios2_fpu_burst_1_upstream_waits_for_read;

  nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register <= NOT nios2_fast_fpu_instruction_master_rdv_fifo_empty_nios2_fpu_burst_1_upstream;
  --local readdatavalid nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream, which is an e_mux
  nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream <= nios2_fpu_burst_1_upstream_readdatavalid_from_sa;
  --byteaddress mux for nios2_fpu_burst_1/upstream, which is an e_mux
  nios2_fpu_burst_1_upstream_byteaddress <= nios2_fast_fpu_instruction_master_address_to_slave (25 DOWNTO 0);
  --master is always granted when requested
  internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream <= internal_nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream;
  --nios2_fast_fpu/instruction_master saved-grant nios2_fpu_burst_1/upstream, which is an e_assign
  nios2_fast_fpu_instruction_master_saved_grant_nios2_fpu_burst_1_upstream <= internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream;
  --allow new arb cycle for nios2_fpu_burst_1/upstream, which is an e_assign
  nios2_fpu_burst_1_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_fpu_burst_1_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_fpu_burst_1_upstream_master_qreq_vector <= std_logic'('1');
  --nios2_fpu_burst_1_upstream_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_1_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_fpu_burst_1_upstream_begins_xfer) = '1'), nios2_fpu_burst_1_upstream_unreg_firsttransfer, nios2_fpu_burst_1_upstream_reg_firsttransfer);
  --nios2_fpu_burst_1_upstream_unreg_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_1_upstream_unreg_firsttransfer <= NOT ((nios2_fpu_burst_1_upstream_slavearbiterlockenable AND nios2_fpu_burst_1_upstream_any_continuerequest));
  --nios2_fpu_burst_1_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_1_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_1_upstream_begins_xfer) = '1' then 
        nios2_fpu_burst_1_upstream_reg_firsttransfer <= nios2_fpu_burst_1_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_1_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_fpu_burst_1_upstream_beginbursttransfer_internal <= nios2_fpu_burst_1_upstream_begins_xfer;
  --nios2_fpu_burst_1_upstream_read assignment, which is an e_mux
  nios2_fpu_burst_1_upstream_read <= internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream AND nios2_fast_fpu_instruction_master_read;
  --nios2_fpu_burst_1_upstream_write assignment, which is an e_mux
  nios2_fpu_burst_1_upstream_write <= std_logic'('0');
  --nios2_fpu_burst_1_upstream_address mux, which is an e_mux
  nios2_fpu_burst_1_upstream_address <= A_EXT (Std_Logic_Vector'(A_SRL(nios2_fast_fpu_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(nios2_fast_fpu_instruction_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 25);
  --d1_nios2_fpu_burst_1_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_fpu_burst_1_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_fpu_burst_1_upstream_end_xfer <= nios2_fpu_burst_1_upstream_end_xfer;
    end if;

  end process;

  --nios2_fpu_burst_1_upstream_waits_for_read in a cycle, which is an e_mux
  nios2_fpu_burst_1_upstream_waits_for_read <= nios2_fpu_burst_1_upstream_in_a_read_cycle AND internal_nios2_fpu_burst_1_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_1_upstream_in_a_read_cycle assignment, which is an e_assign
  nios2_fpu_burst_1_upstream_in_a_read_cycle <= internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream AND nios2_fast_fpu_instruction_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_fpu_burst_1_upstream_in_a_read_cycle;
  --nios2_fpu_burst_1_upstream_waits_for_write in a cycle, which is an e_mux
  nios2_fpu_burst_1_upstream_waits_for_write <= nios2_fpu_burst_1_upstream_in_a_write_cycle AND internal_nios2_fpu_burst_1_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_1_upstream_in_a_write_cycle assignment, which is an e_assign
  nios2_fpu_burst_1_upstream_in_a_write_cycle <= std_logic'('0');
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_fpu_burst_1_upstream_in_a_write_cycle;
  wait_for_nios2_fpu_burst_1_upstream_counter <= std_logic'('0');
  --nios2_fpu_burst_1_upstream_byteenable byte enable port mux, which is an e_mux
  nios2_fpu_burst_1_upstream_byteenable <= A_EXT (-SIGNED(std_logic_vector'("00000000000000000000000000000001")), 2);
  --debugaccess mux, which is an e_mux
  nios2_fpu_burst_1_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream <= internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream;
  --vhdl renameroo for output signals
  nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream <= internal_nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream;
  --vhdl renameroo for output signals
  nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream <= internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream;
  --vhdl renameroo for output signals
  nios2_fpu_burst_1_upstream_waitrequest_from_sa <= internal_nios2_fpu_burst_1_upstream_waitrequest_from_sa;
--synthesis translate_off
    --nios2_fpu_burst_1/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --nios2_fast_fpu/instruction_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line33 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_instruction_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line33, now);
          write(write_line33, string'(": "));
          write(write_line33, string'("nios2_fast_fpu/instruction_master drove 0 on its 'burstcount' port while accessing slave nios2_fpu_burst_1/upstream"));
          write(output, write_line33.all);
          deallocate (write_line33);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_1_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_1_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fpu_burst_1_downstream_granted_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_qualified_request_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_requests_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal nios2_fpu_burst_1_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_1_downstream_latency_counter : OUT STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_1_downstream_readdatavalid : OUT STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_reset_n : OUT STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_waitrequest : OUT STD_LOGIC
              );
end entity nios2_fpu_burst_1_downstream_arbitrator;


architecture europa of nios2_fpu_burst_1_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_fpu_burst_1_downstream_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal internal_nios2_fpu_burst_1_downstream_latency_counter :  STD_LOGIC;
                signal internal_nios2_fpu_burst_1_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_address_last_time :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_1_downstream_burstcount_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fpu_burst_1_downstream_is_granted_some_slave :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_read_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_run :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_write_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_nios2_fpu_burst_1_downstream_latency_counter :  STD_LOGIC;
                signal pre_flush_nios2_fpu_burst_1_downstream_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_1_downstream_qualified_request_sdram_s1 OR NOT nios2_fpu_burst_1_downstream_requests_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_1_downstream_granted_sdram_s1 OR NOT nios2_fpu_burst_1_downstream_qualified_request_sdram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_1_downstream_qualified_request_sdram_s1 OR NOT ((nios2_fpu_burst_1_downstream_read OR nios2_fpu_burst_1_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_1_downstream_read OR nios2_fpu_burst_1_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_1_downstream_qualified_request_sdram_s1 OR NOT ((nios2_fpu_burst_1_downstream_read OR nios2_fpu_burst_1_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_1_downstream_read OR nios2_fpu_burst_1_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_fpu_burst_1_downstream_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_fpu_burst_1_downstream_address_to_slave <= nios2_fpu_burst_1_downstream_address;
  --nios2_fpu_burst_1_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_1_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      nios2_fpu_burst_1_downstream_read_but_no_slave_selected <= (nios2_fpu_burst_1_downstream_read AND nios2_fpu_burst_1_downstream_run) AND NOT nios2_fpu_burst_1_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  nios2_fpu_burst_1_downstream_is_granted_some_slave <= nios2_fpu_burst_1_downstream_granted_sdram_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_nios2_fpu_burst_1_downstream_readdatavalid <= nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  nios2_fpu_burst_1_downstream_readdatavalid <= nios2_fpu_burst_1_downstream_read_but_no_slave_selected OR pre_flush_nios2_fpu_burst_1_downstream_readdatavalid;
  --nios2_fpu_burst_1/downstream readdata mux, which is an e_mux
  nios2_fpu_burst_1_downstream_readdata <= sdram_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_fpu_burst_1_downstream_waitrequest <= NOT nios2_fpu_burst_1_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_nios2_fpu_burst_1_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_nios2_fpu_burst_1_downstream_latency_counter <= p1_nios2_fpu_burst_1_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_nios2_fpu_burst_1_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((nios2_fpu_burst_1_downstream_run AND nios2_fpu_burst_1_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_1_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_1_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --nios2_fpu_burst_1_downstream_reset_n assignment, which is an e_assign
  nios2_fpu_burst_1_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_fpu_burst_1_downstream_address_to_slave <= internal_nios2_fpu_burst_1_downstream_address_to_slave;
  --vhdl renameroo for output signals
  nios2_fpu_burst_1_downstream_latency_counter <= internal_nios2_fpu_burst_1_downstream_latency_counter;
  --vhdl renameroo for output signals
  nios2_fpu_burst_1_downstream_waitrequest <= internal_nios2_fpu_burst_1_downstream_waitrequest;
--synthesis translate_off
    --nios2_fpu_burst_1_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_1_downstream_address_last_time <= std_logic_vector'("0000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_1_downstream_address_last_time <= nios2_fpu_burst_1_downstream_address;
      end if;

    end process;

    --nios2_fpu_burst_1/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_fpu_burst_1_downstream_waitrequest AND ((nios2_fpu_burst_1_downstream_read OR nios2_fpu_burst_1_downstream_write));
      end if;

    end process;

    --nios2_fpu_burst_1_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line34 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_1_downstream_address /= nios2_fpu_burst_1_downstream_address_last_time))))) = '1' then 
          write(write_line34, now);
          write(write_line34, string'(": "));
          write(write_line34, string'("nios2_fpu_burst_1_downstream_address did not heed wait!!!"));
          write(output, write_line34.all);
          deallocate (write_line34);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_1_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_1_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_1_downstream_burstcount_last_time <= nios2_fpu_burst_1_downstream_burstcount;
      end if;

    end process;

    --nios2_fpu_burst_1_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line35 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_1_downstream_burstcount) /= std_logic'(nios2_fpu_burst_1_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line35, now);
          write(write_line35, string'(": "));
          write(write_line35, string'("nios2_fpu_burst_1_downstream_burstcount did not heed wait!!!"));
          write(output, write_line35.all);
          deallocate (write_line35);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_1_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_1_downstream_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_1_downstream_byteenable_last_time <= nios2_fpu_burst_1_downstream_byteenable;
      end if;

    end process;

    --nios2_fpu_burst_1_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line36 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_1_downstream_byteenable /= nios2_fpu_burst_1_downstream_byteenable_last_time))))) = '1' then 
          write(write_line36, now);
          write(write_line36, string'(": "));
          write(write_line36, string'("nios2_fpu_burst_1_downstream_byteenable did not heed wait!!!"));
          write(output, write_line36.all);
          deallocate (write_line36);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_1_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_1_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_1_downstream_read_last_time <= nios2_fpu_burst_1_downstream_read;
      end if;

    end process;

    --nios2_fpu_burst_1_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line37 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_1_downstream_read) /= std_logic'(nios2_fpu_burst_1_downstream_read_last_time)))))) = '1' then 
          write(write_line37, now);
          write(write_line37, string'(": "));
          write(write_line37, string'("nios2_fpu_burst_1_downstream_read did not heed wait!!!"));
          write(output, write_line37.all);
          deallocate (write_line37);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_1_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_1_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_1_downstream_write_last_time <= nios2_fpu_burst_1_downstream_write;
      end if;

    end process;

    --nios2_fpu_burst_1_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line38 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_1_downstream_write) /= std_logic'(nios2_fpu_burst_1_downstream_write_last_time)))))) = '1' then 
          write(write_line38, now);
          write(write_line38, string'(": "));
          write(write_line38, string'("nios2_fpu_burst_1_downstream_write did not heed wait!!!"));
          write(output, write_line38.all);
          deallocate (write_line38);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_1_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_1_downstream_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_1_downstream_writedata_last_time <= nios2_fpu_burst_1_downstream_writedata;
      end if;

    end process;

    --nios2_fpu_burst_1_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line39 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_1_downstream_writedata /= nios2_fpu_burst_1_downstream_writedata_last_time)))) AND nios2_fpu_burst_1_downstream_write)) = '1' then 
          write(write_line39, now);
          write(write_line39, string'(": "));
          write(write_line39, string'("nios2_fpu_burst_1_downstream_writedata did not heed wait!!!"));
          write(output, write_line39.all);
          deallocate (write_line39);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_nios2_fpu_burst_2_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_nios2_fpu_burst_2_upstream_module;


architecture europa of burstcount_fifo_for_nios2_fpu_burst_2_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_3 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_4 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_5 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_6 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_7 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal stage_8 :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_8;
  empty <= NOT(full_0);
  full_9 <= std_logic'('0');
  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic_vector'("00000");
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic_vector'("00000");
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic_vector'("00000");
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic_vector'("00000");
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic_vector'("00000");
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic_vector'("00000");
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("00000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("00000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("00000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 5);
  one_count_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 5);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_2_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_2_upstream_module;


architecture europa of rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_2_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_8;
  empty <= NOT(full_0);
  full_9 <= std_logic'('0');
  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 5);
  one_count_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 5);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_2_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_debugaccess : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_latency_counter : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_2_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_2_upstream_readdatavalid : IN STD_LOGIC;
                 signal nios2_fpu_burst_2_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_nios2_fpu_burst_2_upstream_end_xfer : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream : OUT STD_LOGIC;
                 signal nios2_fpu_burst_2_upstream_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_2_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_2_upstream_byteaddress : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal nios2_fpu_burst_2_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fpu_burst_2_upstream_debugaccess : OUT STD_LOGIC;
                 signal nios2_fpu_burst_2_upstream_read : OUT STD_LOGIC;
                 signal nios2_fpu_burst_2_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_2_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_fpu_burst_2_upstream_write : OUT STD_LOGIC;
                 signal nios2_fpu_burst_2_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity nios2_fpu_burst_2_upstream_arbitrator;


architecture europa of nios2_fpu_burst_2_upstream_arbitrator is
component burstcount_fifo_for_nios2_fpu_burst_2_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_nios2_fpu_burst_2_upstream_module;

component rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_2_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_2_upstream_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_fpu_burst_2_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream :  STD_LOGIC;
                signal internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream :  STD_LOGIC;
                signal internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream :  STD_LOGIC;
                signal internal_nios2_fpu_burst_2_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_nios2_fpu_burst_2_upstream_read :  STD_LOGIC;
                signal internal_nios2_fpu_burst_2_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_nios2_fpu_burst_2_upstream_write :  STD_LOGIC;
                signal module_input12 :  STD_LOGIC;
                signal module_input13 :  STD_LOGIC;
                signal module_input14 :  STD_LOGIC;
                signal module_input15 :  STD_LOGIC;
                signal module_input16 :  STD_LOGIC;
                signal module_input17 :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_arbiterlock :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream_segment_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream_segment_1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_data_master_continuerequest :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_rdv_fifo_empty_nios2_fpu_burst_2_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_rdv_fifo_output_from_nios2_fpu_burst_2_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_saved_grant_nios2_fpu_burst_2_upstream :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_allgrants :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_any_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_arb_counter_enable :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_arb_share_counter :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_begins_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_current_burst :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_end_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_grant_vector :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_in_a_read_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_in_a_write_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_load_fifo :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_master_qreq_vector :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_next_burst_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_reg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_selected_burstcount :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_waits_for_read :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_waits_for_write :  STD_LOGIC;
                signal p0_nios2_fpu_burst_2_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_nios2_fpu_burst_2_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_fpu_burst_2_upstream_end_xfer;
    end if;

  end process;

  nios2_fpu_burst_2_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream);
  --assign nios2_fpu_burst_2_upstream_readdata_from_sa = nios2_fpu_burst_2_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_2_upstream_readdata_from_sa <= nios2_fpu_burst_2_upstream_readdata;
  internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream <= to_std_logic(((Std_Logic_Vector'(nios2_fast_fpu_data_master_address_to_slave(28 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("00000000000000000000000000000")))) AND ((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write));
  --assign nios2_fpu_burst_2_upstream_waitrequest_from_sa = nios2_fpu_burst_2_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_fpu_burst_2_upstream_waitrequest_from_sa <= nios2_fpu_burst_2_upstream_waitrequest;
  --assign nios2_fpu_burst_2_upstream_readdatavalid_from_sa = nios2_fpu_burst_2_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_2_upstream_readdatavalid_from_sa <= nios2_fpu_burst_2_upstream_readdatavalid;
  --nios2_fpu_burst_2_upstream_arb_share_counter set values, which is an e_mux
  nios2_fpu_burst_2_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((nios2_fast_fpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (A_SLL(nios2_fast_fpu_data_master_burstcount,std_logic_vector'("00000000000000000000000000000001")))), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 6);
  --nios2_fpu_burst_2_upstream_non_bursting_master_requests mux, which is an e_mux
  nios2_fpu_burst_2_upstream_non_bursting_master_requests <= std_logic'('0');
  --nios2_fpu_burst_2_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_fpu_burst_2_upstream_any_bursting_master_saved_grant <= nios2_fast_fpu_data_master_saved_grant_nios2_fpu_burst_2_upstream;
  --nios2_fpu_burst_2_upstream_arb_share_counter_next_value assignment, which is an e_assign
  nios2_fpu_burst_2_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_2_upstream_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_2_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_fpu_burst_2_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_2_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 6);
  --nios2_fpu_burst_2_upstream_allgrants all slave grants, which is an e_mux
  nios2_fpu_burst_2_upstream_allgrants <= nios2_fpu_burst_2_upstream_grant_vector;
  --nios2_fpu_burst_2_upstream_end_xfer assignment, which is an e_assign
  nios2_fpu_burst_2_upstream_end_xfer <= NOT ((nios2_fpu_burst_2_upstream_waits_for_read OR nios2_fpu_burst_2_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_fpu_burst_2_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_fpu_burst_2_upstream <= nios2_fpu_burst_2_upstream_end_xfer AND (((NOT nios2_fpu_burst_2_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_fpu_burst_2_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_fpu_burst_2_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_fpu_burst_2_upstream AND nios2_fpu_burst_2_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_2_upstream AND NOT nios2_fpu_burst_2_upstream_non_bursting_master_requests));
  --nios2_fpu_burst_2_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_2_upstream_arb_share_counter <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_2_upstream_arb_counter_enable) = '1' then 
        nios2_fpu_burst_2_upstream_arb_share_counter <= nios2_fpu_burst_2_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_2_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_2_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_fpu_burst_2_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_fpu_burst_2_upstream)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_2_upstream AND NOT nios2_fpu_burst_2_upstream_non_bursting_master_requests)))) = '1' then 
        nios2_fpu_burst_2_upstream_slavearbiterlockenable <= or_reduce(nios2_fpu_burst_2_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --nios2_fast_fpu/data_master nios2_fpu_burst_2/upstream arbiterlock, which is an e_assign
  nios2_fast_fpu_data_master_arbiterlock <= nios2_fpu_burst_2_upstream_slavearbiterlockenable AND nios2_fast_fpu_data_master_continuerequest;
  --nios2_fpu_burst_2_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_fpu_burst_2_upstream_slavearbiterlockenable2 <= or_reduce(nios2_fpu_burst_2_upstream_arb_share_counter_next_value);
  --nios2_fast_fpu/data_master nios2_fpu_burst_2/upstream arbiterlock2, which is an e_assign
  nios2_fast_fpu_data_master_arbiterlock2 <= nios2_fpu_burst_2_upstream_slavearbiterlockenable2 AND nios2_fast_fpu_data_master_continuerequest;
  --nios2_fpu_burst_2_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_fpu_burst_2_upstream_any_continuerequest <= std_logic'('1');
  --nios2_fast_fpu_data_master_continuerequest continued request, which is an e_assign
  nios2_fast_fpu_data_master_continuerequest <= std_logic'('1');
  internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream <= internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream AND NOT ((nios2_fast_fpu_data_master_read AND ((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_data_master_latency_counter))))))) OR (nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register)) OR (nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register)) OR (nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register)))));
  --unique name for nios2_fpu_burst_2_upstream_move_on_to_next_transaction, which is an e_assign
  nios2_fpu_burst_2_upstream_move_on_to_next_transaction <= nios2_fpu_burst_2_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_2_upstream_load_fifo;
  --the currently selected burstcount for nios2_fpu_burst_2_upstream, which is an e_mux
  nios2_fpu_burst_2_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 5);
  --burstcount_fifo_for_nios2_fpu_burst_2_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_nios2_fpu_burst_2_upstream : burstcount_fifo_for_nios2_fpu_burst_2_upstream_module
    port map(
      data_out => nios2_fpu_burst_2_upstream_transaction_burst_count,
      empty => nios2_fpu_burst_2_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input12,
      clk => clk,
      data_in => nios2_fpu_burst_2_upstream_selected_burstcount,
      read => nios2_fpu_burst_2_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input13,
      write => module_input14
    );

  module_input12 <= std_logic'('0');
  module_input13 <= std_logic'('0');
  module_input14 <= ((in_a_read_cycle AND NOT nios2_fpu_burst_2_upstream_waits_for_read) AND nios2_fpu_burst_2_upstream_load_fifo) AND NOT ((nios2_fpu_burst_2_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_2_upstream_burstcount_fifo_empty));

  --nios2_fpu_burst_2_upstream current burst minus one, which is an e_assign
  nios2_fpu_burst_2_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_2_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --what to load in current_burst, for nios2_fpu_burst_2_upstream, which is an e_mux
  nios2_fpu_burst_2_upstream_next_burst_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_2_upstream_waits_for_read)) AND NOT nios2_fpu_burst_2_upstream_load_fifo))) = '1'), (nios2_fpu_burst_2_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_2_upstream_waits_for_read) AND nios2_fpu_burst_2_upstream_this_cycle_is_the_last_burst) AND nios2_fpu_burst_2_upstream_burstcount_fifo_empty))) = '1'), (nios2_fpu_burst_2_upstream_selected_burstcount & A_ToStdLogicVector(std_logic'('0'))), A_WE_StdLogicVector((std_logic'((nios2_fpu_burst_2_upstream_this_cycle_is_the_last_burst)) = '1'), (nios2_fpu_burst_2_upstream_transaction_burst_count & A_ToStdLogicVector(std_logic'('0'))), (std_logic_vector'("0") & (nios2_fpu_burst_2_upstream_current_burst_minus_one))))), 5);
  --the current burst count for nios2_fpu_burst_2_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_2_upstream_current_burst <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((nios2_fpu_burst_2_upstream_readdatavalid_from_sa OR ((NOT nios2_fpu_burst_2_upstream_load_fifo AND ((in_a_read_cycle AND NOT nios2_fpu_burst_2_upstream_waits_for_read)))))) = '1' then 
        nios2_fpu_burst_2_upstream_current_burst <= nios2_fpu_burst_2_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_nios2_fpu_burst_2_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT nios2_fpu_burst_2_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_2_upstream_waits_for_read)) AND nios2_fpu_burst_2_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_2_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_2_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_2_upstream_waits_for_read)) AND NOT nios2_fpu_burst_2_upstream_load_fifo) OR nios2_fpu_burst_2_upstream_this_cycle_is_the_last_burst)) = '1' then 
        nios2_fpu_burst_2_upstream_load_fifo <= p0_nios2_fpu_burst_2_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for nios2_fpu_burst_2_upstream, which is an e_assign
  nios2_fpu_burst_2_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(nios2_fpu_burst_2_upstream_current_burst_minus_one)) AND nios2_fpu_burst_2_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_2_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_2_upstream : rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_2_upstream_module
    port map(
      data_out => nios2_fast_fpu_data_master_rdv_fifo_output_from_nios2_fpu_burst_2_upstream,
      empty => open,
      fifo_contains_ones_n => nios2_fast_fpu_data_master_rdv_fifo_empty_nios2_fpu_burst_2_upstream,
      full => open,
      clear_fifo => module_input15,
      clk => clk,
      data_in => internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream,
      read => nios2_fpu_burst_2_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input16,
      write => module_input17
    );

  module_input15 <= std_logic'('0');
  module_input16 <= std_logic'('0');
  module_input17 <= in_a_read_cycle AND NOT nios2_fpu_burst_2_upstream_waits_for_read;

  nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register <= NOT nios2_fast_fpu_data_master_rdv_fifo_empty_nios2_fpu_burst_2_upstream;
  --local readdatavalid nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream, which is an e_mux
  nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream <= nios2_fpu_burst_2_upstream_readdatavalid_from_sa;
  --nios2_fpu_burst_2_upstream_writedata mux, which is an e_mux
  nios2_fpu_burst_2_upstream_writedata <= nios2_fast_fpu_data_master_dbs_write_16;
  --byteaddress mux for nios2_fpu_burst_2/upstream, which is an e_mux
  nios2_fpu_burst_2_upstream_byteaddress <= nios2_fast_fpu_data_master_address_to_slave (25 DOWNTO 0);
  --master is always granted when requested
  internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream <= internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream;
  --nios2_fast_fpu/data_master saved-grant nios2_fpu_burst_2/upstream, which is an e_assign
  nios2_fast_fpu_data_master_saved_grant_nios2_fpu_burst_2_upstream <= internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream;
  --allow new arb cycle for nios2_fpu_burst_2/upstream, which is an e_assign
  nios2_fpu_burst_2_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_fpu_burst_2_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_fpu_burst_2_upstream_master_qreq_vector <= std_logic'('1');
  --nios2_fpu_burst_2_upstream_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_2_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_fpu_burst_2_upstream_begins_xfer) = '1'), nios2_fpu_burst_2_upstream_unreg_firsttransfer, nios2_fpu_burst_2_upstream_reg_firsttransfer);
  --nios2_fpu_burst_2_upstream_unreg_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_2_upstream_unreg_firsttransfer <= NOT ((nios2_fpu_burst_2_upstream_slavearbiterlockenable AND nios2_fpu_burst_2_upstream_any_continuerequest));
  --nios2_fpu_burst_2_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_2_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_2_upstream_begins_xfer) = '1' then 
        nios2_fpu_burst_2_upstream_reg_firsttransfer <= nios2_fpu_burst_2_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_2_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  nios2_fpu_burst_2_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_nios2_fpu_burst_2_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_2_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_nios2_fpu_burst_2_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_nios2_fpu_burst_2_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_2_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (nios2_fpu_burst_2_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --nios2_fpu_burst_2_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_2_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_2_upstream_begins_xfer) = '1' then 
        nios2_fpu_burst_2_upstream_bbt_burstcounter <= nios2_fpu_burst_2_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_2_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_fpu_burst_2_upstream_beginbursttransfer_internal <= nios2_fpu_burst_2_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_2_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --nios2_fpu_burst_2_upstream_read assignment, which is an e_mux
  internal_nios2_fpu_burst_2_upstream_read <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream AND nios2_fast_fpu_data_master_read;
  --nios2_fpu_burst_2_upstream_write assignment, which is an e_mux
  internal_nios2_fpu_burst_2_upstream_write <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream AND nios2_fast_fpu_data_master_write;
  --nios2_fpu_burst_2_upstream_address mux, which is an e_mux
  nios2_fpu_burst_2_upstream_address <= A_EXT (Std_Logic_Vector'(A_SRL(nios2_fast_fpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(nios2_fast_fpu_data_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 25);
  --d1_nios2_fpu_burst_2_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_fpu_burst_2_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_fpu_burst_2_upstream_end_xfer <= nios2_fpu_burst_2_upstream_end_xfer;
    end if;

  end process;

  --nios2_fpu_burst_2_upstream_waits_for_read in a cycle, which is an e_mux
  nios2_fpu_burst_2_upstream_waits_for_read <= nios2_fpu_burst_2_upstream_in_a_read_cycle AND internal_nios2_fpu_burst_2_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_2_upstream_in_a_read_cycle assignment, which is an e_assign
  nios2_fpu_burst_2_upstream_in_a_read_cycle <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream AND nios2_fast_fpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_fpu_burst_2_upstream_in_a_read_cycle;
  --nios2_fpu_burst_2_upstream_waits_for_write in a cycle, which is an e_mux
  nios2_fpu_burst_2_upstream_waits_for_write <= nios2_fpu_burst_2_upstream_in_a_write_cycle AND internal_nios2_fpu_burst_2_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_2_upstream_in_a_write_cycle assignment, which is an e_assign
  nios2_fpu_burst_2_upstream_in_a_write_cycle <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream AND nios2_fast_fpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_fpu_burst_2_upstream_in_a_write_cycle;
  wait_for_nios2_fpu_burst_2_upstream_counter <= std_logic'('0');
  --nios2_fpu_burst_2_upstream_byteenable byte enable port mux, which is an e_mux
  nios2_fpu_burst_2_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (internal_nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  (nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream_segment_1(1), nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream_segment_1(0), nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream_segment_0(1), nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream_segment_0(0)) <= nios2_fast_fpu_data_master_byteenable;
  internal_nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_data_master_dbs_address(1)))) = std_logic_vector'("00000000000000000000000000000000"))), nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream_segment_0, nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream_segment_1);
  --burstcount mux, which is an e_mux
  internal_nios2_fpu_burst_2_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  nios2_fpu_burst_2_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream <= internal_nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream;
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream;
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream <= internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream;
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream <= internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream;
  --vhdl renameroo for output signals
  nios2_fpu_burst_2_upstream_burstcount <= internal_nios2_fpu_burst_2_upstream_burstcount;
  --vhdl renameroo for output signals
  nios2_fpu_burst_2_upstream_read <= internal_nios2_fpu_burst_2_upstream_read;
  --vhdl renameroo for output signals
  nios2_fpu_burst_2_upstream_waitrequest_from_sa <= internal_nios2_fpu_burst_2_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  nios2_fpu_burst_2_upstream_write <= internal_nios2_fpu_burst_2_upstream_write;
--synthesis translate_off
    --nios2_fpu_burst_2/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --nios2_fast_fpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line40 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line40, now);
          write(write_line40, string'(": "));
          write(write_line40, string'("nios2_fast_fpu/data_master drove 0 on its 'burstcount' port while accessing slave nios2_fpu_burst_2/upstream"));
          write(output, write_line40.all);
          deallocate (write_line40);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_2_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_2_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fpu_burst_2_downstream_granted_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_qualified_request_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_requests_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal nios2_fpu_burst_2_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_2_downstream_latency_counter : OUT STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_2_downstream_readdatavalid : OUT STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_reset_n : OUT STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_waitrequest : OUT STD_LOGIC
              );
end entity nios2_fpu_burst_2_downstream_arbitrator;


architecture europa of nios2_fpu_burst_2_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_fpu_burst_2_downstream_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal internal_nios2_fpu_burst_2_downstream_latency_counter :  STD_LOGIC;
                signal internal_nios2_fpu_burst_2_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_address_last_time :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_2_downstream_burstcount_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fpu_burst_2_downstream_is_granted_some_slave :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_read_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_run :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_write_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_nios2_fpu_burst_2_downstream_latency_counter :  STD_LOGIC;
                signal pre_flush_nios2_fpu_burst_2_downstream_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_2_downstream_qualified_request_sdram_s1 OR NOT nios2_fpu_burst_2_downstream_requests_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_2_downstream_granted_sdram_s1 OR NOT nios2_fpu_burst_2_downstream_qualified_request_sdram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_2_downstream_qualified_request_sdram_s1 OR NOT ((nios2_fpu_burst_2_downstream_read OR nios2_fpu_burst_2_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_2_downstream_read OR nios2_fpu_burst_2_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_2_downstream_qualified_request_sdram_s1 OR NOT ((nios2_fpu_burst_2_downstream_read OR nios2_fpu_burst_2_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_2_downstream_read OR nios2_fpu_burst_2_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_fpu_burst_2_downstream_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_fpu_burst_2_downstream_address_to_slave <= nios2_fpu_burst_2_downstream_address;
  --nios2_fpu_burst_2_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_2_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      nios2_fpu_burst_2_downstream_read_but_no_slave_selected <= (nios2_fpu_burst_2_downstream_read AND nios2_fpu_burst_2_downstream_run) AND NOT nios2_fpu_burst_2_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  nios2_fpu_burst_2_downstream_is_granted_some_slave <= nios2_fpu_burst_2_downstream_granted_sdram_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_nios2_fpu_burst_2_downstream_readdatavalid <= nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  nios2_fpu_burst_2_downstream_readdatavalid <= nios2_fpu_burst_2_downstream_read_but_no_slave_selected OR pre_flush_nios2_fpu_burst_2_downstream_readdatavalid;
  --nios2_fpu_burst_2/downstream readdata mux, which is an e_mux
  nios2_fpu_burst_2_downstream_readdata <= sdram_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_fpu_burst_2_downstream_waitrequest <= NOT nios2_fpu_burst_2_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_nios2_fpu_burst_2_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_nios2_fpu_burst_2_downstream_latency_counter <= p1_nios2_fpu_burst_2_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_nios2_fpu_burst_2_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((nios2_fpu_burst_2_downstream_run AND nios2_fpu_burst_2_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_2_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_2_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --nios2_fpu_burst_2_downstream_reset_n assignment, which is an e_assign
  nios2_fpu_burst_2_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_fpu_burst_2_downstream_address_to_slave <= internal_nios2_fpu_burst_2_downstream_address_to_slave;
  --vhdl renameroo for output signals
  nios2_fpu_burst_2_downstream_latency_counter <= internal_nios2_fpu_burst_2_downstream_latency_counter;
  --vhdl renameroo for output signals
  nios2_fpu_burst_2_downstream_waitrequest <= internal_nios2_fpu_burst_2_downstream_waitrequest;
--synthesis translate_off
    --nios2_fpu_burst_2_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_2_downstream_address_last_time <= std_logic_vector'("0000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_2_downstream_address_last_time <= nios2_fpu_burst_2_downstream_address;
      end if;

    end process;

    --nios2_fpu_burst_2/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_fpu_burst_2_downstream_waitrequest AND ((nios2_fpu_burst_2_downstream_read OR nios2_fpu_burst_2_downstream_write));
      end if;

    end process;

    --nios2_fpu_burst_2_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line41 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_2_downstream_address /= nios2_fpu_burst_2_downstream_address_last_time))))) = '1' then 
          write(write_line41, now);
          write(write_line41, string'(": "));
          write(write_line41, string'("nios2_fpu_burst_2_downstream_address did not heed wait!!!"));
          write(output, write_line41.all);
          deallocate (write_line41);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_2_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_2_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_2_downstream_burstcount_last_time <= nios2_fpu_burst_2_downstream_burstcount;
      end if;

    end process;

    --nios2_fpu_burst_2_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line42 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_2_downstream_burstcount) /= std_logic'(nios2_fpu_burst_2_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line42, now);
          write(write_line42, string'(": "));
          write(write_line42, string'("nios2_fpu_burst_2_downstream_burstcount did not heed wait!!!"));
          write(output, write_line42.all);
          deallocate (write_line42);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_2_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_2_downstream_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_2_downstream_byteenable_last_time <= nios2_fpu_burst_2_downstream_byteenable;
      end if;

    end process;

    --nios2_fpu_burst_2_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line43 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_2_downstream_byteenable /= nios2_fpu_burst_2_downstream_byteenable_last_time))))) = '1' then 
          write(write_line43, now);
          write(write_line43, string'(": "));
          write(write_line43, string'("nios2_fpu_burst_2_downstream_byteenable did not heed wait!!!"));
          write(output, write_line43.all);
          deallocate (write_line43);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_2_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_2_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_2_downstream_read_last_time <= nios2_fpu_burst_2_downstream_read;
      end if;

    end process;

    --nios2_fpu_burst_2_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line44 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_2_downstream_read) /= std_logic'(nios2_fpu_burst_2_downstream_read_last_time)))))) = '1' then 
          write(write_line44, now);
          write(write_line44, string'(": "));
          write(write_line44, string'("nios2_fpu_burst_2_downstream_read did not heed wait!!!"));
          write(output, write_line44.all);
          deallocate (write_line44);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_2_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_2_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_2_downstream_write_last_time <= nios2_fpu_burst_2_downstream_write;
      end if;

    end process;

    --nios2_fpu_burst_2_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line45 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_2_downstream_write) /= std_logic'(nios2_fpu_burst_2_downstream_write_last_time)))))) = '1' then 
          write(write_line45, now);
          write(write_line45, string'(": "));
          write(write_line45, string'("nios2_fpu_burst_2_downstream_write did not heed wait!!!"));
          write(output, write_line45.all);
          deallocate (write_line45);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_2_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_2_downstream_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_2_downstream_writedata_last_time <= nios2_fpu_burst_2_downstream_writedata;
      end if;

    end process;

    --nios2_fpu_burst_2_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line46 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_2_downstream_writedata /= nios2_fpu_burst_2_downstream_writedata_last_time)))) AND nios2_fpu_burst_2_downstream_write)) = '1' then 
          write(write_line46, now);
          write(write_line46, string'(": "));
          write(write_line46, string'("nios2_fpu_burst_2_downstream_writedata did not heed wait!!!"));
          write(output, write_line46.all);
          deallocate (write_line46);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_nios2_fpu_burst_3_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_nios2_fpu_burst_3_upstream_module;


architecture europa of burstcount_fifo_for_nios2_fpu_burst_3_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_3 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_4 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_5 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_6 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_7 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_8 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_8;
  empty <= NOT(full_0);
  full_9 <= std_logic'('0');
  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic_vector'("000");
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic_vector'("000");
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic_vector'("000");
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic_vector'("000");
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic_vector'("000");
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic_vector'("000");
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 5);
  one_count_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 5);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_spu_m1_to_nios2_fpu_burst_3_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_spu_m1_to_nios2_fpu_burst_3_upstream_module;


architecture europa of rdv_fifo_for_spu_m1_to_nios2_fpu_burst_3_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_8;
  empty <= NOT(full_0);
  full_9 <= std_logic'('0');
  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 5);
  one_count_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 5);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_3_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_3_upstream_readdatavalid : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal spu_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal spu_m1_burstcount : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal spu_m1_latency_counter : IN STD_LOGIC;
                 signal spu_m1_read : IN STD_LOGIC;

              -- outputs:
                 signal d1_nios2_fpu_burst_3_upstream_end_xfer : OUT STD_LOGIC;
                 signal nios2_fpu_burst_3_upstream_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_3_upstream_burstcount : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_fpu_burst_3_upstream_byteaddress : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal nios2_fpu_burst_3_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fpu_burst_3_upstream_debugaccess : OUT STD_LOGIC;
                 signal nios2_fpu_burst_3_upstream_read : OUT STD_LOGIC;
                 signal nios2_fpu_burst_3_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_3_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_fpu_burst_3_upstream_write : OUT STD_LOGIC;
                 signal spu_m1_granted_nios2_fpu_burst_3_upstream : OUT STD_LOGIC;
                 signal spu_m1_qualified_request_nios2_fpu_burst_3_upstream : OUT STD_LOGIC;
                 signal spu_m1_read_data_valid_nios2_fpu_burst_3_upstream : OUT STD_LOGIC;
                 signal spu_m1_read_data_valid_nios2_fpu_burst_3_upstream_shift_register : OUT STD_LOGIC;
                 signal spu_m1_requests_nios2_fpu_burst_3_upstream : OUT STD_LOGIC
              );
end entity nios2_fpu_burst_3_upstream_arbitrator;


architecture europa of nios2_fpu_burst_3_upstream_arbitrator is
component burstcount_fifo_for_nios2_fpu_burst_3_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_nios2_fpu_burst_3_upstream_module;

component rdv_fifo_for_spu_m1_to_nios2_fpu_burst_3_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_spu_m1_to_nios2_fpu_burst_3_upstream_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_fpu_burst_3_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_fpu_burst_3_upstream_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_nios2_fpu_burst_3_upstream_read :  STD_LOGIC;
                signal internal_nios2_fpu_burst_3_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_nios2_fpu_burst_3_upstream_write :  STD_LOGIC;
                signal internal_spu_m1_granted_nios2_fpu_burst_3_upstream :  STD_LOGIC;
                signal internal_spu_m1_qualified_request_nios2_fpu_burst_3_upstream :  STD_LOGIC;
                signal internal_spu_m1_requests_nios2_fpu_burst_3_upstream :  STD_LOGIC;
                signal module_input18 :  STD_LOGIC;
                signal module_input19 :  STD_LOGIC;
                signal module_input20 :  STD_LOGIC;
                signal module_input21 :  STD_LOGIC;
                signal module_input22 :  STD_LOGIC;
                signal module_input23 :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_allgrants :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_any_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_arb_counter_enable :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_begins_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_current_burst :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_end_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_grant_vector :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_in_a_read_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_in_a_write_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_load_fifo :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_master_qreq_vector :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_next_burst_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_reg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_selected_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_waits_for_read :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_waits_for_write :  STD_LOGIC;
                signal p0_nios2_fpu_burst_3_upstream_load_fifo :  STD_LOGIC;
                signal spu_m1_arbiterlock :  STD_LOGIC;
                signal spu_m1_arbiterlock2 :  STD_LOGIC;
                signal spu_m1_continuerequest :  STD_LOGIC;
                signal spu_m1_rdv_fifo_empty_nios2_fpu_burst_3_upstream :  STD_LOGIC;
                signal spu_m1_rdv_fifo_output_from_nios2_fpu_burst_3_upstream :  STD_LOGIC;
                signal spu_m1_saved_grant_nios2_fpu_burst_3_upstream :  STD_LOGIC;
                signal wait_for_nios2_fpu_burst_3_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_fpu_burst_3_upstream_end_xfer;
    end if;

  end process;

  nios2_fpu_burst_3_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_spu_m1_qualified_request_nios2_fpu_burst_3_upstream);
  --assign nios2_fpu_burst_3_upstream_readdata_from_sa = nios2_fpu_burst_3_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_3_upstream_readdata_from_sa <= nios2_fpu_burst_3_upstream_readdata;
  internal_spu_m1_requests_nios2_fpu_burst_3_upstream <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((spu_m1_read)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(spu_m1_read)))));
  --assign nios2_fpu_burst_3_upstream_waitrequest_from_sa = nios2_fpu_burst_3_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_fpu_burst_3_upstream_waitrequest_from_sa <= nios2_fpu_burst_3_upstream_waitrequest;
  --assign nios2_fpu_burst_3_upstream_readdatavalid_from_sa = nios2_fpu_burst_3_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_3_upstream_readdatavalid_from_sa <= nios2_fpu_burst_3_upstream_readdatavalid;
  --nios2_fpu_burst_3_upstream_arb_share_counter set values, which is an e_mux
  nios2_fpu_burst_3_upstream_arb_share_set_values <= std_logic_vector'("001");
  --nios2_fpu_burst_3_upstream_non_bursting_master_requests mux, which is an e_mux
  nios2_fpu_burst_3_upstream_non_bursting_master_requests <= std_logic'('0');
  --nios2_fpu_burst_3_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_fpu_burst_3_upstream_any_bursting_master_saved_grant <= spu_m1_saved_grant_nios2_fpu_burst_3_upstream;
  --nios2_fpu_burst_3_upstream_arb_share_counter_next_value assignment, which is an e_assign
  nios2_fpu_burst_3_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_3_upstream_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (nios2_fpu_burst_3_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_fpu_burst_3_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (nios2_fpu_burst_3_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --nios2_fpu_burst_3_upstream_allgrants all slave grants, which is an e_mux
  nios2_fpu_burst_3_upstream_allgrants <= nios2_fpu_burst_3_upstream_grant_vector;
  --nios2_fpu_burst_3_upstream_end_xfer assignment, which is an e_assign
  nios2_fpu_burst_3_upstream_end_xfer <= NOT ((nios2_fpu_burst_3_upstream_waits_for_read OR nios2_fpu_burst_3_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_fpu_burst_3_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_fpu_burst_3_upstream <= nios2_fpu_burst_3_upstream_end_xfer AND (((NOT nios2_fpu_burst_3_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_fpu_burst_3_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_fpu_burst_3_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_fpu_burst_3_upstream AND nios2_fpu_burst_3_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_3_upstream AND NOT nios2_fpu_burst_3_upstream_non_bursting_master_requests));
  --nios2_fpu_burst_3_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_3_upstream_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_3_upstream_arb_counter_enable) = '1' then 
        nios2_fpu_burst_3_upstream_arb_share_counter <= nios2_fpu_burst_3_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_3_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_3_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_fpu_burst_3_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_fpu_burst_3_upstream)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_3_upstream AND NOT nios2_fpu_burst_3_upstream_non_bursting_master_requests)))) = '1' then 
        nios2_fpu_burst_3_upstream_slavearbiterlockenable <= or_reduce(nios2_fpu_burst_3_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --spu/m1 nios2_fpu_burst_3/upstream arbiterlock, which is an e_assign
  spu_m1_arbiterlock <= nios2_fpu_burst_3_upstream_slavearbiterlockenable AND spu_m1_continuerequest;
  --nios2_fpu_burst_3_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_fpu_burst_3_upstream_slavearbiterlockenable2 <= or_reduce(nios2_fpu_burst_3_upstream_arb_share_counter_next_value);
  --spu/m1 nios2_fpu_burst_3/upstream arbiterlock2, which is an e_assign
  spu_m1_arbiterlock2 <= nios2_fpu_burst_3_upstream_slavearbiterlockenable2 AND spu_m1_continuerequest;
  --nios2_fpu_burst_3_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_fpu_burst_3_upstream_any_continuerequest <= std_logic'('1');
  --spu_m1_continuerequest continued request, which is an e_assign
  spu_m1_continuerequest <= std_logic'('1');
  internal_spu_m1_qualified_request_nios2_fpu_burst_3_upstream <= internal_spu_m1_requests_nios2_fpu_burst_3_upstream AND NOT ((spu_m1_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(spu_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(spu_m1_latency_counter))))))))));
  --unique name for nios2_fpu_burst_3_upstream_move_on_to_next_transaction, which is an e_assign
  nios2_fpu_burst_3_upstream_move_on_to_next_transaction <= nios2_fpu_burst_3_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_3_upstream_load_fifo;
  --the currently selected burstcount for nios2_fpu_burst_3_upstream, which is an e_mux
  nios2_fpu_burst_3_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_spu_m1_granted_nios2_fpu_burst_3_upstream)) = '1'), (std_logic_vector'("00000000000000000000000000000") & (spu_m1_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 3);
  --burstcount_fifo_for_nios2_fpu_burst_3_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_nios2_fpu_burst_3_upstream : burstcount_fifo_for_nios2_fpu_burst_3_upstream_module
    port map(
      data_out => nios2_fpu_burst_3_upstream_transaction_burst_count,
      empty => nios2_fpu_burst_3_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input18,
      clk => clk,
      data_in => nios2_fpu_burst_3_upstream_selected_burstcount,
      read => nios2_fpu_burst_3_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input19,
      write => module_input20
    );

  module_input18 <= std_logic'('0');
  module_input19 <= std_logic'('0');
  module_input20 <= ((in_a_read_cycle AND NOT nios2_fpu_burst_3_upstream_waits_for_read) AND nios2_fpu_burst_3_upstream_load_fifo) AND NOT ((nios2_fpu_burst_3_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_3_upstream_burstcount_fifo_empty));

  --nios2_fpu_burst_3_upstream current burst minus one, which is an e_assign
  nios2_fpu_burst_3_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (nios2_fpu_burst_3_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --what to load in current_burst, for nios2_fpu_burst_3_upstream, which is an e_mux
  nios2_fpu_burst_3_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_3_upstream_waits_for_read)) AND NOT nios2_fpu_burst_3_upstream_load_fifo))) = '1'), nios2_fpu_burst_3_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_3_upstream_waits_for_read) AND nios2_fpu_burst_3_upstream_this_cycle_is_the_last_burst) AND nios2_fpu_burst_3_upstream_burstcount_fifo_empty))) = '1'), nios2_fpu_burst_3_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((nios2_fpu_burst_3_upstream_this_cycle_is_the_last_burst)) = '1'), nios2_fpu_burst_3_upstream_transaction_burst_count, nios2_fpu_burst_3_upstream_current_burst_minus_one)));
  --the current burst count for nios2_fpu_burst_3_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_3_upstream_current_burst <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((nios2_fpu_burst_3_upstream_readdatavalid_from_sa OR ((NOT nios2_fpu_burst_3_upstream_load_fifo AND ((in_a_read_cycle AND NOT nios2_fpu_burst_3_upstream_waits_for_read)))))) = '1' then 
        nios2_fpu_burst_3_upstream_current_burst <= nios2_fpu_burst_3_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_nios2_fpu_burst_3_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT nios2_fpu_burst_3_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_3_upstream_waits_for_read)) AND nios2_fpu_burst_3_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_3_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_3_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_3_upstream_waits_for_read)) AND NOT nios2_fpu_burst_3_upstream_load_fifo) OR nios2_fpu_burst_3_upstream_this_cycle_is_the_last_burst)) = '1' then 
        nios2_fpu_burst_3_upstream_load_fifo <= p0_nios2_fpu_burst_3_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for nios2_fpu_burst_3_upstream, which is an e_assign
  nios2_fpu_burst_3_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(nios2_fpu_burst_3_upstream_current_burst_minus_one)) AND nios2_fpu_burst_3_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_spu_m1_to_nios2_fpu_burst_3_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_spu_m1_to_nios2_fpu_burst_3_upstream : rdv_fifo_for_spu_m1_to_nios2_fpu_burst_3_upstream_module
    port map(
      data_out => spu_m1_rdv_fifo_output_from_nios2_fpu_burst_3_upstream,
      empty => open,
      fifo_contains_ones_n => spu_m1_rdv_fifo_empty_nios2_fpu_burst_3_upstream,
      full => open,
      clear_fifo => module_input21,
      clk => clk,
      data_in => internal_spu_m1_granted_nios2_fpu_burst_3_upstream,
      read => nios2_fpu_burst_3_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input22,
      write => module_input23
    );

  module_input21 <= std_logic'('0');
  module_input22 <= std_logic'('0');
  module_input23 <= in_a_read_cycle AND NOT nios2_fpu_burst_3_upstream_waits_for_read;

  spu_m1_read_data_valid_nios2_fpu_burst_3_upstream_shift_register <= NOT spu_m1_rdv_fifo_empty_nios2_fpu_burst_3_upstream;
  --local readdatavalid spu_m1_read_data_valid_nios2_fpu_burst_3_upstream, which is an e_mux
  spu_m1_read_data_valid_nios2_fpu_burst_3_upstream <= nios2_fpu_burst_3_upstream_readdatavalid_from_sa;
  --byteaddress mux for nios2_fpu_burst_3/upstream, which is an e_mux
  nios2_fpu_burst_3_upstream_byteaddress <= std_logic_vector'("0") & (spu_m1_address_to_slave);
  --master is always granted when requested
  internal_spu_m1_granted_nios2_fpu_burst_3_upstream <= internal_spu_m1_qualified_request_nios2_fpu_burst_3_upstream;
  --spu/m1 saved-grant nios2_fpu_burst_3/upstream, which is an e_assign
  spu_m1_saved_grant_nios2_fpu_burst_3_upstream <= internal_spu_m1_requests_nios2_fpu_burst_3_upstream;
  --allow new arb cycle for nios2_fpu_burst_3/upstream, which is an e_assign
  nios2_fpu_burst_3_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_fpu_burst_3_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_fpu_burst_3_upstream_master_qreq_vector <= std_logic'('1');
  --nios2_fpu_burst_3_upstream_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_3_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_fpu_burst_3_upstream_begins_xfer) = '1'), nios2_fpu_burst_3_upstream_unreg_firsttransfer, nios2_fpu_burst_3_upstream_reg_firsttransfer);
  --nios2_fpu_burst_3_upstream_unreg_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_3_upstream_unreg_firsttransfer <= NOT ((nios2_fpu_burst_3_upstream_slavearbiterlockenable AND nios2_fpu_burst_3_upstream_any_continuerequest));
  --nios2_fpu_burst_3_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_3_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_3_upstream_begins_xfer) = '1' then 
        nios2_fpu_burst_3_upstream_reg_firsttransfer <= nios2_fpu_burst_3_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_3_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  nios2_fpu_burst_3_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_nios2_fpu_burst_3_upstream_write) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (nios2_fpu_burst_3_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (internal_nios2_fpu_burst_3_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_nios2_fpu_burst_3_upstream_read) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (nios2_fpu_burst_3_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("0000000000000000000000000000000") & (nios2_fpu_burst_3_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 2);
  --nios2_fpu_burst_3_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_3_upstream_bbt_burstcounter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_3_upstream_begins_xfer) = '1' then 
        nios2_fpu_burst_3_upstream_bbt_burstcounter <= nios2_fpu_burst_3_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_3_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_fpu_burst_3_upstream_beginbursttransfer_internal <= nios2_fpu_burst_3_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (nios2_fpu_burst_3_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --nios2_fpu_burst_3_upstream_read assignment, which is an e_mux
  internal_nios2_fpu_burst_3_upstream_read <= internal_spu_m1_granted_nios2_fpu_burst_3_upstream AND spu_m1_read;
  --nios2_fpu_burst_3_upstream_write assignment, which is an e_mux
  internal_nios2_fpu_burst_3_upstream_write <= std_logic'('0');
  --nios2_fpu_burst_3_upstream_address mux, which is an e_mux
  nios2_fpu_burst_3_upstream_address <= spu_m1_address_to_slave;
  --d1_nios2_fpu_burst_3_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_fpu_burst_3_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_fpu_burst_3_upstream_end_xfer <= nios2_fpu_burst_3_upstream_end_xfer;
    end if;

  end process;

  --nios2_fpu_burst_3_upstream_waits_for_read in a cycle, which is an e_mux
  nios2_fpu_burst_3_upstream_waits_for_read <= nios2_fpu_burst_3_upstream_in_a_read_cycle AND internal_nios2_fpu_burst_3_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_3_upstream_in_a_read_cycle assignment, which is an e_assign
  nios2_fpu_burst_3_upstream_in_a_read_cycle <= internal_spu_m1_granted_nios2_fpu_burst_3_upstream AND spu_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_fpu_burst_3_upstream_in_a_read_cycle;
  --nios2_fpu_burst_3_upstream_waits_for_write in a cycle, which is an e_mux
  nios2_fpu_burst_3_upstream_waits_for_write <= nios2_fpu_burst_3_upstream_in_a_write_cycle AND internal_nios2_fpu_burst_3_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_3_upstream_in_a_write_cycle assignment, which is an e_assign
  nios2_fpu_burst_3_upstream_in_a_write_cycle <= std_logic'('0');
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_fpu_burst_3_upstream_in_a_write_cycle;
  wait_for_nios2_fpu_burst_3_upstream_counter <= std_logic'('0');
  --nios2_fpu_burst_3_upstream_byteenable byte enable port mux, which is an e_mux
  nios2_fpu_burst_3_upstream_byteenable <= A_EXT (-SIGNED(std_logic_vector'("00000000000000000000000000000001")), 2);
  --burstcount mux, which is an e_mux
  internal_nios2_fpu_burst_3_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_spu_m1_granted_nios2_fpu_burst_3_upstream)) = '1'), (std_logic_vector'("00000000000000000000000000000") & (spu_m1_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 3);
  --debugaccess mux, which is an e_mux
  nios2_fpu_burst_3_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_fpu_burst_3_upstream_burstcount <= internal_nios2_fpu_burst_3_upstream_burstcount;
  --vhdl renameroo for output signals
  nios2_fpu_burst_3_upstream_read <= internal_nios2_fpu_burst_3_upstream_read;
  --vhdl renameroo for output signals
  nios2_fpu_burst_3_upstream_waitrequest_from_sa <= internal_nios2_fpu_burst_3_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  nios2_fpu_burst_3_upstream_write <= internal_nios2_fpu_burst_3_upstream_write;
  --vhdl renameroo for output signals
  spu_m1_granted_nios2_fpu_burst_3_upstream <= internal_spu_m1_granted_nios2_fpu_burst_3_upstream;
  --vhdl renameroo for output signals
  spu_m1_qualified_request_nios2_fpu_burst_3_upstream <= internal_spu_m1_qualified_request_nios2_fpu_burst_3_upstream;
  --vhdl renameroo for output signals
  spu_m1_requests_nios2_fpu_burst_3_upstream <= internal_spu_m1_requests_nios2_fpu_burst_3_upstream;
--synthesis translate_off
    --nios2_fpu_burst_3/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --spu/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line47 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_spu_m1_requests_nios2_fpu_burst_3_upstream AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (spu_m1_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line47, now);
          write(write_line47, string'(": "));
          write(write_line47, string'("spu/m1 drove 0 on its 'burstcount' port while accessing slave nios2_fpu_burst_3/upstream"));
          write(output, write_line47.all);
          deallocate (write_line47);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_3_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_3_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fpu_burst_3_downstream_granted_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_qualified_request_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_requests_sdram_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal nios2_fpu_burst_3_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_3_downstream_latency_counter : OUT STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_3_downstream_readdatavalid : OUT STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_reset_n : OUT STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_waitrequest : OUT STD_LOGIC
              );
end entity nios2_fpu_burst_3_downstream_arbitrator;


architecture europa of nios2_fpu_burst_3_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_fpu_burst_3_downstream_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal internal_nios2_fpu_burst_3_downstream_latency_counter :  STD_LOGIC;
                signal internal_nios2_fpu_burst_3_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_address_last_time :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_3_downstream_burstcount_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fpu_burst_3_downstream_is_granted_some_slave :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_read_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_run :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_write_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_nios2_fpu_burst_3_downstream_latency_counter :  STD_LOGIC;
                signal pre_flush_nios2_fpu_burst_3_downstream_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_3_downstream_qualified_request_sdram_s1 OR NOT nios2_fpu_burst_3_downstream_requests_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_3_downstream_granted_sdram_s1 OR NOT nios2_fpu_burst_3_downstream_qualified_request_sdram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_3_downstream_qualified_request_sdram_s1 OR NOT ((nios2_fpu_burst_3_downstream_read OR nios2_fpu_burst_3_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_3_downstream_read OR nios2_fpu_burst_3_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_3_downstream_qualified_request_sdram_s1 OR NOT ((nios2_fpu_burst_3_downstream_read OR nios2_fpu_burst_3_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_3_downstream_read OR nios2_fpu_burst_3_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_fpu_burst_3_downstream_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_fpu_burst_3_downstream_address_to_slave <= nios2_fpu_burst_3_downstream_address;
  --nios2_fpu_burst_3_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_3_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      nios2_fpu_burst_3_downstream_read_but_no_slave_selected <= (nios2_fpu_burst_3_downstream_read AND nios2_fpu_burst_3_downstream_run) AND NOT nios2_fpu_burst_3_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  nios2_fpu_burst_3_downstream_is_granted_some_slave <= nios2_fpu_burst_3_downstream_granted_sdram_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_nios2_fpu_burst_3_downstream_readdatavalid <= nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  nios2_fpu_burst_3_downstream_readdatavalid <= nios2_fpu_burst_3_downstream_read_but_no_slave_selected OR pre_flush_nios2_fpu_burst_3_downstream_readdatavalid;
  --nios2_fpu_burst_3/downstream readdata mux, which is an e_mux
  nios2_fpu_burst_3_downstream_readdata <= sdram_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_fpu_burst_3_downstream_waitrequest <= NOT nios2_fpu_burst_3_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_nios2_fpu_burst_3_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_nios2_fpu_burst_3_downstream_latency_counter <= p1_nios2_fpu_burst_3_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_nios2_fpu_burst_3_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((nios2_fpu_burst_3_downstream_run AND nios2_fpu_burst_3_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_3_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_3_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --nios2_fpu_burst_3_downstream_reset_n assignment, which is an e_assign
  nios2_fpu_burst_3_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_fpu_burst_3_downstream_address_to_slave <= internal_nios2_fpu_burst_3_downstream_address_to_slave;
  --vhdl renameroo for output signals
  nios2_fpu_burst_3_downstream_latency_counter <= internal_nios2_fpu_burst_3_downstream_latency_counter;
  --vhdl renameroo for output signals
  nios2_fpu_burst_3_downstream_waitrequest <= internal_nios2_fpu_burst_3_downstream_waitrequest;
--synthesis translate_off
    --nios2_fpu_burst_3_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_3_downstream_address_last_time <= std_logic_vector'("0000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_3_downstream_address_last_time <= nios2_fpu_burst_3_downstream_address;
      end if;

    end process;

    --nios2_fpu_burst_3/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_fpu_burst_3_downstream_waitrequest AND ((nios2_fpu_burst_3_downstream_read OR nios2_fpu_burst_3_downstream_write));
      end if;

    end process;

    --nios2_fpu_burst_3_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line48 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_3_downstream_address /= nios2_fpu_burst_3_downstream_address_last_time))))) = '1' then 
          write(write_line48, now);
          write(write_line48, string'(": "));
          write(write_line48, string'("nios2_fpu_burst_3_downstream_address did not heed wait!!!"));
          write(output, write_line48.all);
          deallocate (write_line48);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_3_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_3_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_3_downstream_burstcount_last_time <= nios2_fpu_burst_3_downstream_burstcount;
      end if;

    end process;

    --nios2_fpu_burst_3_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line49 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_3_downstream_burstcount) /= std_logic'(nios2_fpu_burst_3_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line49, now);
          write(write_line49, string'(": "));
          write(write_line49, string'("nios2_fpu_burst_3_downstream_burstcount did not heed wait!!!"));
          write(output, write_line49.all);
          deallocate (write_line49);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_3_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_3_downstream_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_3_downstream_byteenable_last_time <= nios2_fpu_burst_3_downstream_byteenable;
      end if;

    end process;

    --nios2_fpu_burst_3_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line50 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_3_downstream_byteenable /= nios2_fpu_burst_3_downstream_byteenable_last_time))))) = '1' then 
          write(write_line50, now);
          write(write_line50, string'(": "));
          write(write_line50, string'("nios2_fpu_burst_3_downstream_byteenable did not heed wait!!!"));
          write(output, write_line50.all);
          deallocate (write_line50);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_3_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_3_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_3_downstream_read_last_time <= nios2_fpu_burst_3_downstream_read;
      end if;

    end process;

    --nios2_fpu_burst_3_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line51 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_3_downstream_read) /= std_logic'(nios2_fpu_burst_3_downstream_read_last_time)))))) = '1' then 
          write(write_line51, now);
          write(write_line51, string'(": "));
          write(write_line51, string'("nios2_fpu_burst_3_downstream_read did not heed wait!!!"));
          write(output, write_line51.all);
          deallocate (write_line51);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_3_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_3_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_3_downstream_write_last_time <= nios2_fpu_burst_3_downstream_write;
      end if;

    end process;

    --nios2_fpu_burst_3_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line52 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_3_downstream_write) /= std_logic'(nios2_fpu_burst_3_downstream_write_last_time)))))) = '1' then 
          write(write_line52, now);
          write(write_line52, string'(": "));
          write(write_line52, string'("nios2_fpu_burst_3_downstream_write did not heed wait!!!"));
          write(output, write_line52.all);
          deallocate (write_line52);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_3_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_3_downstream_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_3_downstream_writedata_last_time <= nios2_fpu_burst_3_downstream_writedata;
      end if;

    end process;

    --nios2_fpu_burst_3_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line53 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_3_downstream_writedata /= nios2_fpu_burst_3_downstream_writedata_last_time)))) AND nios2_fpu_burst_3_downstream_write)) = '1' then 
          write(write_line53, now);
          write(write_line53, string'(": "));
          write(write_line53, string'("nios2_fpu_burst_3_downstream_writedata did not heed wait!!!"));
          write(output, write_line53.all);
          deallocate (write_line53);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_nios2_fpu_burst_4_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_nios2_fpu_burst_4_upstream_module;


architecture europa of burstcount_fifo_for_nios2_fpu_burst_4_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_4_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_4_upstream_module;


architecture europa of rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_4_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_4_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal nios2_fast_fpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fast_fpu_instruction_master_latency_counter : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_4_upstream_readdatavalid : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_nios2_fpu_burst_4_upstream_end_xfer : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream : OUT STD_LOGIC;
                 signal nios2_fpu_burst_4_upstream_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal nios2_fpu_burst_4_upstream_byteaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_burst_4_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_4_upstream_debugaccess : OUT STD_LOGIC;
                 signal nios2_fpu_burst_4_upstream_read : OUT STD_LOGIC;
                 signal nios2_fpu_burst_4_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_4_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_fpu_burst_4_upstream_write : OUT STD_LOGIC
              );
end entity nios2_fpu_burst_4_upstream_arbitrator;


architecture europa of nios2_fpu_burst_4_upstream_arbitrator is
component burstcount_fifo_for_nios2_fpu_burst_4_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_nios2_fpu_burst_4_upstream_module;

component rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_4_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_4_upstream_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_fpu_burst_4_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream :  STD_LOGIC;
                signal internal_nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream :  STD_LOGIC;
                signal internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream :  STD_LOGIC;
                signal internal_nios2_fpu_burst_4_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal module_input24 :  STD_LOGIC;
                signal module_input25 :  STD_LOGIC;
                signal module_input26 :  STD_LOGIC;
                signal module_input27 :  STD_LOGIC;
                signal module_input28 :  STD_LOGIC;
                signal module_input29 :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_continuerequest :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_rdv_fifo_empty_nios2_fpu_burst_4_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_rdv_fifo_output_from_nios2_fpu_burst_4_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_saved_grant_nios2_fpu_burst_4_upstream :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_allgrants :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_any_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_arb_counter_enable :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_arb_share_counter :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_4_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_4_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_4_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_begins_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_4_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_4_upstream_end_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_grant_vector :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_in_a_read_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_in_a_write_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_load_fifo :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_master_qreq_vector :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_4_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_reg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_4_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_4_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_waits_for_read :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_waits_for_write :  STD_LOGIC;
                signal p0_nios2_fpu_burst_4_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_nios2_fpu_burst_4_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_fpu_burst_4_upstream_end_xfer;
    end if;

  end process;

  nios2_fpu_burst_4_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream);
  --assign nios2_fpu_burst_4_upstream_readdatavalid_from_sa = nios2_fpu_burst_4_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_4_upstream_readdatavalid_from_sa <= nios2_fpu_burst_4_upstream_readdatavalid;
  --assign nios2_fpu_burst_4_upstream_readdata_from_sa = nios2_fpu_burst_4_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_4_upstream_readdata_from_sa <= nios2_fpu_burst_4_upstream_readdata;
  internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream <= ((to_std_logic(((Std_Logic_Vector'(nios2_fast_fpu_instruction_master_address_to_slave(27 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("1111111111110000100000000000")))) AND (nios2_fast_fpu_instruction_master_read))) AND nios2_fast_fpu_instruction_master_read;
  --assign nios2_fpu_burst_4_upstream_waitrequest_from_sa = nios2_fpu_burst_4_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_fpu_burst_4_upstream_waitrequest_from_sa <= nios2_fpu_burst_4_upstream_waitrequest;
  --nios2_fpu_burst_4_upstream_arb_share_counter set values, which is an e_mux
  nios2_fpu_burst_4_upstream_arb_share_set_values <= std_logic_vector'("000001");
  --nios2_fpu_burst_4_upstream_non_bursting_master_requests mux, which is an e_mux
  nios2_fpu_burst_4_upstream_non_bursting_master_requests <= std_logic'('0');
  --nios2_fpu_burst_4_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_fpu_burst_4_upstream_any_bursting_master_saved_grant <= nios2_fast_fpu_instruction_master_saved_grant_nios2_fpu_burst_4_upstream;
  --nios2_fpu_burst_4_upstream_arb_share_counter_next_value assignment, which is an e_assign
  nios2_fpu_burst_4_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_4_upstream_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_4_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_fpu_burst_4_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_4_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 6);
  --nios2_fpu_burst_4_upstream_allgrants all slave grants, which is an e_mux
  nios2_fpu_burst_4_upstream_allgrants <= nios2_fpu_burst_4_upstream_grant_vector;
  --nios2_fpu_burst_4_upstream_end_xfer assignment, which is an e_assign
  nios2_fpu_burst_4_upstream_end_xfer <= NOT ((nios2_fpu_burst_4_upstream_waits_for_read OR nios2_fpu_burst_4_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_fpu_burst_4_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_fpu_burst_4_upstream <= nios2_fpu_burst_4_upstream_end_xfer AND (((NOT nios2_fpu_burst_4_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_fpu_burst_4_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_fpu_burst_4_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_fpu_burst_4_upstream AND nios2_fpu_burst_4_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_4_upstream AND NOT nios2_fpu_burst_4_upstream_non_bursting_master_requests));
  --nios2_fpu_burst_4_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_4_upstream_arb_share_counter <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_4_upstream_arb_counter_enable) = '1' then 
        nios2_fpu_burst_4_upstream_arb_share_counter <= nios2_fpu_burst_4_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_4_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_4_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_fpu_burst_4_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_fpu_burst_4_upstream)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_4_upstream AND NOT nios2_fpu_burst_4_upstream_non_bursting_master_requests)))) = '1' then 
        nios2_fpu_burst_4_upstream_slavearbiterlockenable <= or_reduce(nios2_fpu_burst_4_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --nios2_fast_fpu/instruction_master nios2_fpu_burst_4/upstream arbiterlock, which is an e_assign
  nios2_fast_fpu_instruction_master_arbiterlock <= nios2_fpu_burst_4_upstream_slavearbiterlockenable AND nios2_fast_fpu_instruction_master_continuerequest;
  --nios2_fpu_burst_4_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_fpu_burst_4_upstream_slavearbiterlockenable2 <= or_reduce(nios2_fpu_burst_4_upstream_arb_share_counter_next_value);
  --nios2_fast_fpu/instruction_master nios2_fpu_burst_4/upstream arbiterlock2, which is an e_assign
  nios2_fast_fpu_instruction_master_arbiterlock2 <= nios2_fpu_burst_4_upstream_slavearbiterlockenable2 AND nios2_fast_fpu_instruction_master_continuerequest;
  --nios2_fpu_burst_4_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_fpu_burst_4_upstream_any_continuerequest <= std_logic'('1');
  --nios2_fast_fpu_instruction_master_continuerequest continued request, which is an e_assign
  nios2_fast_fpu_instruction_master_continuerequest <= std_logic'('1');
  internal_nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream <= internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream AND NOT ((nios2_fast_fpu_instruction_master_read AND (((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_instruction_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_instruction_master_latency_counter))))))) OR (nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register)) OR (nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register)))));
  --unique name for nios2_fpu_burst_4_upstream_move_on_to_next_transaction, which is an e_assign
  nios2_fpu_burst_4_upstream_move_on_to_next_transaction <= nios2_fpu_burst_4_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_4_upstream_load_fifo;
  --the currently selected burstcount for nios2_fpu_burst_4_upstream, which is an e_mux
  nios2_fpu_burst_4_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_instruction_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_nios2_fpu_burst_4_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_nios2_fpu_burst_4_upstream : burstcount_fifo_for_nios2_fpu_burst_4_upstream_module
    port map(
      data_out => nios2_fpu_burst_4_upstream_transaction_burst_count,
      empty => nios2_fpu_burst_4_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input24,
      clk => clk,
      data_in => nios2_fpu_burst_4_upstream_selected_burstcount,
      read => nios2_fpu_burst_4_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input25,
      write => module_input26
    );

  module_input24 <= std_logic'('0');
  module_input25 <= std_logic'('0');
  module_input26 <= ((in_a_read_cycle AND NOT nios2_fpu_burst_4_upstream_waits_for_read) AND nios2_fpu_burst_4_upstream_load_fifo) AND NOT ((nios2_fpu_burst_4_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_4_upstream_burstcount_fifo_empty));

  --nios2_fpu_burst_4_upstream current burst minus one, which is an e_assign
  nios2_fpu_burst_4_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_4_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for nios2_fpu_burst_4_upstream, which is an e_mux
  nios2_fpu_burst_4_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_4_upstream_waits_for_read)) AND NOT nios2_fpu_burst_4_upstream_load_fifo))) = '1'), nios2_fpu_burst_4_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_4_upstream_waits_for_read) AND nios2_fpu_burst_4_upstream_this_cycle_is_the_last_burst) AND nios2_fpu_burst_4_upstream_burstcount_fifo_empty))) = '1'), nios2_fpu_burst_4_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((nios2_fpu_burst_4_upstream_this_cycle_is_the_last_burst)) = '1'), nios2_fpu_burst_4_upstream_transaction_burst_count, nios2_fpu_burst_4_upstream_current_burst_minus_one)));
  --the current burst count for nios2_fpu_burst_4_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_4_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((nios2_fpu_burst_4_upstream_readdatavalid_from_sa OR ((NOT nios2_fpu_burst_4_upstream_load_fifo AND ((in_a_read_cycle AND NOT nios2_fpu_burst_4_upstream_waits_for_read)))))) = '1' then 
        nios2_fpu_burst_4_upstream_current_burst <= nios2_fpu_burst_4_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_nios2_fpu_burst_4_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT nios2_fpu_burst_4_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_4_upstream_waits_for_read)) AND nios2_fpu_burst_4_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_4_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_4_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_4_upstream_waits_for_read)) AND NOT nios2_fpu_burst_4_upstream_load_fifo) OR nios2_fpu_burst_4_upstream_this_cycle_is_the_last_burst)) = '1' then 
        nios2_fpu_burst_4_upstream_load_fifo <= p0_nios2_fpu_burst_4_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for nios2_fpu_burst_4_upstream, which is an e_assign
  nios2_fpu_burst_4_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(nios2_fpu_burst_4_upstream_current_burst_minus_one)) AND nios2_fpu_burst_4_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_4_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_4_upstream : rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_4_upstream_module
    port map(
      data_out => nios2_fast_fpu_instruction_master_rdv_fifo_output_from_nios2_fpu_burst_4_upstream,
      empty => open,
      fifo_contains_ones_n => nios2_fast_fpu_instruction_master_rdv_fifo_empty_nios2_fpu_burst_4_upstream,
      full => open,
      clear_fifo => module_input27,
      clk => clk,
      data_in => internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream,
      read => nios2_fpu_burst_4_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input28,
      write => module_input29
    );

  module_input27 <= std_logic'('0');
  module_input28 <= std_logic'('0');
  module_input29 <= in_a_read_cycle AND NOT nios2_fpu_burst_4_upstream_waits_for_read;

  nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register <= NOT nios2_fast_fpu_instruction_master_rdv_fifo_empty_nios2_fpu_burst_4_upstream;
  --local readdatavalid nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream, which is an e_mux
  nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream <= nios2_fpu_burst_4_upstream_readdatavalid_from_sa;
  --byteaddress mux for nios2_fpu_burst_4/upstream, which is an e_mux
  nios2_fpu_burst_4_upstream_byteaddress <= nios2_fast_fpu_instruction_master_address_to_slave (12 DOWNTO 0);
  --master is always granted when requested
  internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream <= internal_nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream;
  --nios2_fast_fpu/instruction_master saved-grant nios2_fpu_burst_4/upstream, which is an e_assign
  nios2_fast_fpu_instruction_master_saved_grant_nios2_fpu_burst_4_upstream <= internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream;
  --allow new arb cycle for nios2_fpu_burst_4/upstream, which is an e_assign
  nios2_fpu_burst_4_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_fpu_burst_4_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_fpu_burst_4_upstream_master_qreq_vector <= std_logic'('1');
  --nios2_fpu_burst_4_upstream_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_4_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_fpu_burst_4_upstream_begins_xfer) = '1'), nios2_fpu_burst_4_upstream_unreg_firsttransfer, nios2_fpu_burst_4_upstream_reg_firsttransfer);
  --nios2_fpu_burst_4_upstream_unreg_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_4_upstream_unreg_firsttransfer <= NOT ((nios2_fpu_burst_4_upstream_slavearbiterlockenable AND nios2_fpu_burst_4_upstream_any_continuerequest));
  --nios2_fpu_burst_4_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_4_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_4_upstream_begins_xfer) = '1' then 
        nios2_fpu_burst_4_upstream_reg_firsttransfer <= nios2_fpu_burst_4_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_4_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_fpu_burst_4_upstream_beginbursttransfer_internal <= nios2_fpu_burst_4_upstream_begins_xfer;
  --nios2_fpu_burst_4_upstream_read assignment, which is an e_mux
  nios2_fpu_burst_4_upstream_read <= internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream AND nios2_fast_fpu_instruction_master_read;
  --nios2_fpu_burst_4_upstream_write assignment, which is an e_mux
  nios2_fpu_burst_4_upstream_write <= std_logic'('0');
  --nios2_fpu_burst_4_upstream_address mux, which is an e_mux
  nios2_fpu_burst_4_upstream_address <= nios2_fast_fpu_instruction_master_address_to_slave (10 DOWNTO 0);
  --d1_nios2_fpu_burst_4_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_fpu_burst_4_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_fpu_burst_4_upstream_end_xfer <= nios2_fpu_burst_4_upstream_end_xfer;
    end if;

  end process;

  --nios2_fpu_burst_4_upstream_waits_for_read in a cycle, which is an e_mux
  nios2_fpu_burst_4_upstream_waits_for_read <= nios2_fpu_burst_4_upstream_in_a_read_cycle AND internal_nios2_fpu_burst_4_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_4_upstream_in_a_read_cycle assignment, which is an e_assign
  nios2_fpu_burst_4_upstream_in_a_read_cycle <= internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream AND nios2_fast_fpu_instruction_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_fpu_burst_4_upstream_in_a_read_cycle;
  --nios2_fpu_burst_4_upstream_waits_for_write in a cycle, which is an e_mux
  nios2_fpu_burst_4_upstream_waits_for_write <= nios2_fpu_burst_4_upstream_in_a_write_cycle AND internal_nios2_fpu_burst_4_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_4_upstream_in_a_write_cycle assignment, which is an e_assign
  nios2_fpu_burst_4_upstream_in_a_write_cycle <= std_logic'('0');
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_fpu_burst_4_upstream_in_a_write_cycle;
  wait_for_nios2_fpu_burst_4_upstream_counter <= std_logic'('0');
  --nios2_fpu_burst_4_upstream_byteenable byte enable port mux, which is an e_mux
  nios2_fpu_burst_4_upstream_byteenable <= A_EXT (-SIGNED(std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  nios2_fpu_burst_4_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream <= internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream;
  --vhdl renameroo for output signals
  nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream <= internal_nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream;
  --vhdl renameroo for output signals
  nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream <= internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream;
  --vhdl renameroo for output signals
  nios2_fpu_burst_4_upstream_waitrequest_from_sa <= internal_nios2_fpu_burst_4_upstream_waitrequest_from_sa;
--synthesis translate_off
    --nios2_fpu_burst_4/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --nios2_fast_fpu/instruction_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line54 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_instruction_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line54, now);
          write(write_line54, string'(": "));
          write(write_line54, string'("nios2_fast_fpu/instruction_master drove 0 on its 'burstcount' port while accessing slave nios2_fpu_burst_4/upstream"));
          write(output, write_line54.all);
          deallocate (write_line54);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_4_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_nios2_fast_fpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal nios2_fast_fpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_4_downstream_address : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal nios2_fpu_burst_4_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_fpu_burst_4_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal nios2_fpu_burst_4_downstream_latency_counter : OUT STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_4_downstream_readdatavalid : OUT STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_reset_n : OUT STD_LOGIC;
                 signal nios2_fpu_burst_4_downstream_waitrequest : OUT STD_LOGIC
              );
end entity nios2_fpu_burst_4_downstream_arbitrator;


architecture europa of nios2_fpu_burst_4_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_fpu_burst_4_downstream_address_to_slave :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal internal_nios2_fpu_burst_4_downstream_latency_counter :  STD_LOGIC;
                signal internal_nios2_fpu_burst_4_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_address_last_time :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_4_downstream_burstcount_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_4_downstream_is_granted_some_slave :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_read_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_run :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_write_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_nios2_fpu_burst_4_downstream_latency_counter :  STD_LOGIC;
                signal pre_flush_nios2_fpu_burst_4_downstream_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module OR NOT nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module OR NOT nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module OR NOT nios2_fpu_burst_4_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_nios2_fast_fpu_jtag_debug_module_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_4_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module OR NOT nios2_fpu_burst_4_downstream_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_4_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_fpu_burst_4_downstream_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_fpu_burst_4_downstream_address_to_slave <= nios2_fpu_burst_4_downstream_address;
  --nios2_fpu_burst_4_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_4_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      nios2_fpu_burst_4_downstream_read_but_no_slave_selected <= (nios2_fpu_burst_4_downstream_read AND nios2_fpu_burst_4_downstream_run) AND NOT nios2_fpu_burst_4_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  nios2_fpu_burst_4_downstream_is_granted_some_slave <= nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_nios2_fpu_burst_4_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  nios2_fpu_burst_4_downstream_readdatavalid <= (nios2_fpu_burst_4_downstream_read_but_no_slave_selected OR pre_flush_nios2_fpu_burst_4_downstream_readdatavalid) OR nios2_fpu_burst_4_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module;
  --nios2_fpu_burst_4/downstream readdata mux, which is an e_mux
  nios2_fpu_burst_4_downstream_readdata <= nios2_fast_fpu_jtag_debug_module_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_fpu_burst_4_downstream_waitrequest <= NOT nios2_fpu_burst_4_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_nios2_fpu_burst_4_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_nios2_fpu_burst_4_downstream_latency_counter <= p1_nios2_fpu_burst_4_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_nios2_fpu_burst_4_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((nios2_fpu_burst_4_downstream_run AND nios2_fpu_burst_4_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_4_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_4_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --nios2_fpu_burst_4_downstream_reset_n assignment, which is an e_assign
  nios2_fpu_burst_4_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_fpu_burst_4_downstream_address_to_slave <= internal_nios2_fpu_burst_4_downstream_address_to_slave;
  --vhdl renameroo for output signals
  nios2_fpu_burst_4_downstream_latency_counter <= internal_nios2_fpu_burst_4_downstream_latency_counter;
  --vhdl renameroo for output signals
  nios2_fpu_burst_4_downstream_waitrequest <= internal_nios2_fpu_burst_4_downstream_waitrequest;
--synthesis translate_off
    --nios2_fpu_burst_4_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_4_downstream_address_last_time <= std_logic_vector'("00000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_4_downstream_address_last_time <= nios2_fpu_burst_4_downstream_address;
      end if;

    end process;

    --nios2_fpu_burst_4/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_fpu_burst_4_downstream_waitrequest AND ((nios2_fpu_burst_4_downstream_read OR nios2_fpu_burst_4_downstream_write));
      end if;

    end process;

    --nios2_fpu_burst_4_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line55 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_4_downstream_address /= nios2_fpu_burst_4_downstream_address_last_time))))) = '1' then 
          write(write_line55, now);
          write(write_line55, string'(": "));
          write(write_line55, string'("nios2_fpu_burst_4_downstream_address did not heed wait!!!"));
          write(output, write_line55.all);
          deallocate (write_line55);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_4_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_4_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_4_downstream_burstcount_last_time <= nios2_fpu_burst_4_downstream_burstcount;
      end if;

    end process;

    --nios2_fpu_burst_4_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line56 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_4_downstream_burstcount) /= std_logic'(nios2_fpu_burst_4_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line56, now);
          write(write_line56, string'(": "));
          write(write_line56, string'("nios2_fpu_burst_4_downstream_burstcount did not heed wait!!!"));
          write(output, write_line56.all);
          deallocate (write_line56);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_4_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_4_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_4_downstream_byteenable_last_time <= nios2_fpu_burst_4_downstream_byteenable;
      end if;

    end process;

    --nios2_fpu_burst_4_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line57 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_4_downstream_byteenable /= nios2_fpu_burst_4_downstream_byteenable_last_time))))) = '1' then 
          write(write_line57, now);
          write(write_line57, string'(": "));
          write(write_line57, string'("nios2_fpu_burst_4_downstream_byteenable did not heed wait!!!"));
          write(output, write_line57.all);
          deallocate (write_line57);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_4_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_4_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_4_downstream_read_last_time <= nios2_fpu_burst_4_downstream_read;
      end if;

    end process;

    --nios2_fpu_burst_4_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line58 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_4_downstream_read) /= std_logic'(nios2_fpu_burst_4_downstream_read_last_time)))))) = '1' then 
          write(write_line58, now);
          write(write_line58, string'(": "));
          write(write_line58, string'("nios2_fpu_burst_4_downstream_read did not heed wait!!!"));
          write(output, write_line58.all);
          deallocate (write_line58);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_4_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_4_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_4_downstream_write_last_time <= nios2_fpu_burst_4_downstream_write;
      end if;

    end process;

    --nios2_fpu_burst_4_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line59 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_4_downstream_write) /= std_logic'(nios2_fpu_burst_4_downstream_write_last_time)))))) = '1' then 
          write(write_line59, now);
          write(write_line59, string'(": "));
          write(write_line59, string'("nios2_fpu_burst_4_downstream_write did not heed wait!!!"));
          write(output, write_line59.all);
          deallocate (write_line59);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_4_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_4_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_4_downstream_writedata_last_time <= nios2_fpu_burst_4_downstream_writedata;
      end if;

    end process;

    --nios2_fpu_burst_4_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line60 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_4_downstream_writedata /= nios2_fpu_burst_4_downstream_writedata_last_time)))) AND nios2_fpu_burst_4_downstream_write)) = '1' then 
          write(write_line60, now);
          write(write_line60, string'(": "));
          write(write_line60, string'("nios2_fpu_burst_4_downstream_writedata did not heed wait!!!"));
          write(output, write_line60.all);
          deallocate (write_line60);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_nios2_fpu_burst_5_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_nios2_fpu_burst_5_upstream_module;


architecture europa of burstcount_fifo_for_nios2_fpu_burst_5_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_5_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_5_upstream_module;


architecture europa of rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_5_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_1;
  empty <= NOT(full_0);
  full_2 <= std_logic'('0');
  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_0))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_5_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_debugaccess : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_latency_counter : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_write : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_5_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_5_upstream_readdatavalid : IN STD_LOGIC;
                 signal nios2_fpu_burst_5_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_nios2_fpu_burst_5_upstream_end_xfer : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream : OUT STD_LOGIC;
                 signal nios2_fpu_burst_5_upstream_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal nios2_fpu_burst_5_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_5_upstream_byteaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_burst_5_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_5_upstream_debugaccess : OUT STD_LOGIC;
                 signal nios2_fpu_burst_5_upstream_read : OUT STD_LOGIC;
                 signal nios2_fpu_burst_5_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_5_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_fpu_burst_5_upstream_write : OUT STD_LOGIC;
                 signal nios2_fpu_burst_5_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity nios2_fpu_burst_5_upstream_arbitrator;


architecture europa of nios2_fpu_burst_5_upstream_arbitrator is
component burstcount_fifo_for_nios2_fpu_burst_5_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_nios2_fpu_burst_5_upstream_module;

component rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_5_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_5_upstream_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_fpu_burst_5_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream :  STD_LOGIC;
                signal internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream :  STD_LOGIC;
                signal internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream :  STD_LOGIC;
                signal internal_nios2_fpu_burst_5_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_nios2_fpu_burst_5_upstream_read :  STD_LOGIC;
                signal internal_nios2_fpu_burst_5_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_nios2_fpu_burst_5_upstream_write :  STD_LOGIC;
                signal module_input30 :  STD_LOGIC;
                signal module_input31 :  STD_LOGIC;
                signal module_input32 :  STD_LOGIC;
                signal module_input33 :  STD_LOGIC;
                signal module_input34 :  STD_LOGIC;
                signal module_input35 :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_arbiterlock :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_continuerequest :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_rdv_fifo_empty_nios2_fpu_burst_5_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_rdv_fifo_output_from_nios2_fpu_burst_5_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_saved_grant_nios2_fpu_burst_5_upstream :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_allgrants :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_any_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_arb_counter_enable :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_arb_share_counter :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_begins_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_end_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_grant_vector :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_in_a_read_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_in_a_write_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_load_fifo :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_master_qreq_vector :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_reg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_waits_for_read :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_waits_for_write :  STD_LOGIC;
                signal p0_nios2_fpu_burst_5_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_nios2_fpu_burst_5_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_fpu_burst_5_upstream_end_xfer;
    end if;

  end process;

  nios2_fpu_burst_5_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream);
  --assign nios2_fpu_burst_5_upstream_readdatavalid_from_sa = nios2_fpu_burst_5_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_5_upstream_readdatavalid_from_sa <= nios2_fpu_burst_5_upstream_readdatavalid;
  --assign nios2_fpu_burst_5_upstream_readdata_from_sa = nios2_fpu_burst_5_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_5_upstream_readdata_from_sa <= nios2_fpu_burst_5_upstream_readdata;
  internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream <= to_std_logic(((Std_Logic_Vector'(nios2_fast_fpu_data_master_address_to_slave(28 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("01111111111110000100000000000")))) AND ((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write));
  --assign nios2_fpu_burst_5_upstream_waitrequest_from_sa = nios2_fpu_burst_5_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_fpu_burst_5_upstream_waitrequest_from_sa <= nios2_fpu_burst_5_upstream_waitrequest;
  --nios2_fpu_burst_5_upstream_arb_share_counter set values, which is an e_mux
  nios2_fpu_burst_5_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((nios2_fast_fpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 6);
  --nios2_fpu_burst_5_upstream_non_bursting_master_requests mux, which is an e_mux
  nios2_fpu_burst_5_upstream_non_bursting_master_requests <= std_logic'('0');
  --nios2_fpu_burst_5_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_fpu_burst_5_upstream_any_bursting_master_saved_grant <= nios2_fast_fpu_data_master_saved_grant_nios2_fpu_burst_5_upstream;
  --nios2_fpu_burst_5_upstream_arb_share_counter_next_value assignment, which is an e_assign
  nios2_fpu_burst_5_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_5_upstream_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_5_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_fpu_burst_5_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_5_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 6);
  --nios2_fpu_burst_5_upstream_allgrants all slave grants, which is an e_mux
  nios2_fpu_burst_5_upstream_allgrants <= nios2_fpu_burst_5_upstream_grant_vector;
  --nios2_fpu_burst_5_upstream_end_xfer assignment, which is an e_assign
  nios2_fpu_burst_5_upstream_end_xfer <= NOT ((nios2_fpu_burst_5_upstream_waits_for_read OR nios2_fpu_burst_5_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_fpu_burst_5_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_fpu_burst_5_upstream <= nios2_fpu_burst_5_upstream_end_xfer AND (((NOT nios2_fpu_burst_5_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_fpu_burst_5_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_fpu_burst_5_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_fpu_burst_5_upstream AND nios2_fpu_burst_5_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_5_upstream AND NOT nios2_fpu_burst_5_upstream_non_bursting_master_requests));
  --nios2_fpu_burst_5_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_5_upstream_arb_share_counter <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_5_upstream_arb_counter_enable) = '1' then 
        nios2_fpu_burst_5_upstream_arb_share_counter <= nios2_fpu_burst_5_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_5_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_5_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_fpu_burst_5_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_fpu_burst_5_upstream)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_5_upstream AND NOT nios2_fpu_burst_5_upstream_non_bursting_master_requests)))) = '1' then 
        nios2_fpu_burst_5_upstream_slavearbiterlockenable <= or_reduce(nios2_fpu_burst_5_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --nios2_fast_fpu/data_master nios2_fpu_burst_5/upstream arbiterlock, which is an e_assign
  nios2_fast_fpu_data_master_arbiterlock <= nios2_fpu_burst_5_upstream_slavearbiterlockenable AND nios2_fast_fpu_data_master_continuerequest;
  --nios2_fpu_burst_5_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_fpu_burst_5_upstream_slavearbiterlockenable2 <= or_reduce(nios2_fpu_burst_5_upstream_arb_share_counter_next_value);
  --nios2_fast_fpu/data_master nios2_fpu_burst_5/upstream arbiterlock2, which is an e_assign
  nios2_fast_fpu_data_master_arbiterlock2 <= nios2_fpu_burst_5_upstream_slavearbiterlockenable2 AND nios2_fast_fpu_data_master_continuerequest;
  --nios2_fpu_burst_5_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_fpu_burst_5_upstream_any_continuerequest <= std_logic'('1');
  --nios2_fast_fpu_data_master_continuerequest continued request, which is an e_assign
  nios2_fast_fpu_data_master_continuerequest <= std_logic'('1');
  internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream <= internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream AND NOT ((nios2_fast_fpu_data_master_read AND ((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_data_master_latency_counter))))))) OR (nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register)) OR (nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register)) OR (nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register)))));
  --unique name for nios2_fpu_burst_5_upstream_move_on_to_next_transaction, which is an e_assign
  nios2_fpu_burst_5_upstream_move_on_to_next_transaction <= nios2_fpu_burst_5_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_5_upstream_load_fifo;
  --the currently selected burstcount for nios2_fpu_burst_5_upstream, which is an e_mux
  nios2_fpu_burst_5_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_nios2_fpu_burst_5_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_nios2_fpu_burst_5_upstream : burstcount_fifo_for_nios2_fpu_burst_5_upstream_module
    port map(
      data_out => nios2_fpu_burst_5_upstream_transaction_burst_count,
      empty => nios2_fpu_burst_5_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input30,
      clk => clk,
      data_in => nios2_fpu_burst_5_upstream_selected_burstcount,
      read => nios2_fpu_burst_5_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input31,
      write => module_input32
    );

  module_input30 <= std_logic'('0');
  module_input31 <= std_logic'('0');
  module_input32 <= ((in_a_read_cycle AND NOT nios2_fpu_burst_5_upstream_waits_for_read) AND nios2_fpu_burst_5_upstream_load_fifo) AND NOT ((nios2_fpu_burst_5_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_5_upstream_burstcount_fifo_empty));

  --nios2_fpu_burst_5_upstream current burst minus one, which is an e_assign
  nios2_fpu_burst_5_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_5_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for nios2_fpu_burst_5_upstream, which is an e_mux
  nios2_fpu_burst_5_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_5_upstream_waits_for_read)) AND NOT nios2_fpu_burst_5_upstream_load_fifo))) = '1'), nios2_fpu_burst_5_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_5_upstream_waits_for_read) AND nios2_fpu_burst_5_upstream_this_cycle_is_the_last_burst) AND nios2_fpu_burst_5_upstream_burstcount_fifo_empty))) = '1'), nios2_fpu_burst_5_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((nios2_fpu_burst_5_upstream_this_cycle_is_the_last_burst)) = '1'), nios2_fpu_burst_5_upstream_transaction_burst_count, nios2_fpu_burst_5_upstream_current_burst_minus_one)));
  --the current burst count for nios2_fpu_burst_5_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_5_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((nios2_fpu_burst_5_upstream_readdatavalid_from_sa OR ((NOT nios2_fpu_burst_5_upstream_load_fifo AND ((in_a_read_cycle AND NOT nios2_fpu_burst_5_upstream_waits_for_read)))))) = '1' then 
        nios2_fpu_burst_5_upstream_current_burst <= nios2_fpu_burst_5_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_nios2_fpu_burst_5_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT nios2_fpu_burst_5_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_5_upstream_waits_for_read)) AND nios2_fpu_burst_5_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_5_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_5_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_5_upstream_waits_for_read)) AND NOT nios2_fpu_burst_5_upstream_load_fifo) OR nios2_fpu_burst_5_upstream_this_cycle_is_the_last_burst)) = '1' then 
        nios2_fpu_burst_5_upstream_load_fifo <= p0_nios2_fpu_burst_5_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for nios2_fpu_burst_5_upstream, which is an e_assign
  nios2_fpu_burst_5_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(nios2_fpu_burst_5_upstream_current_burst_minus_one)) AND nios2_fpu_burst_5_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_5_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_5_upstream : rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_5_upstream_module
    port map(
      data_out => nios2_fast_fpu_data_master_rdv_fifo_output_from_nios2_fpu_burst_5_upstream,
      empty => open,
      fifo_contains_ones_n => nios2_fast_fpu_data_master_rdv_fifo_empty_nios2_fpu_burst_5_upstream,
      full => open,
      clear_fifo => module_input33,
      clk => clk,
      data_in => internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream,
      read => nios2_fpu_burst_5_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input34,
      write => module_input35
    );

  module_input33 <= std_logic'('0');
  module_input34 <= std_logic'('0');
  module_input35 <= in_a_read_cycle AND NOT nios2_fpu_burst_5_upstream_waits_for_read;

  nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register <= NOT nios2_fast_fpu_data_master_rdv_fifo_empty_nios2_fpu_burst_5_upstream;
  --local readdatavalid nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream, which is an e_mux
  nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream <= nios2_fpu_burst_5_upstream_readdatavalid_from_sa;
  --nios2_fpu_burst_5_upstream_writedata mux, which is an e_mux
  nios2_fpu_burst_5_upstream_writedata <= nios2_fast_fpu_data_master_writedata;
  --byteaddress mux for nios2_fpu_burst_5/upstream, which is an e_mux
  nios2_fpu_burst_5_upstream_byteaddress <= nios2_fast_fpu_data_master_address_to_slave (12 DOWNTO 0);
  --master is always granted when requested
  internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream <= internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream;
  --nios2_fast_fpu/data_master saved-grant nios2_fpu_burst_5/upstream, which is an e_assign
  nios2_fast_fpu_data_master_saved_grant_nios2_fpu_burst_5_upstream <= internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream;
  --allow new arb cycle for nios2_fpu_burst_5/upstream, which is an e_assign
  nios2_fpu_burst_5_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_fpu_burst_5_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_fpu_burst_5_upstream_master_qreq_vector <= std_logic'('1');
  --nios2_fpu_burst_5_upstream_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_5_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_fpu_burst_5_upstream_begins_xfer) = '1'), nios2_fpu_burst_5_upstream_unreg_firsttransfer, nios2_fpu_burst_5_upstream_reg_firsttransfer);
  --nios2_fpu_burst_5_upstream_unreg_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_5_upstream_unreg_firsttransfer <= NOT ((nios2_fpu_burst_5_upstream_slavearbiterlockenable AND nios2_fpu_burst_5_upstream_any_continuerequest));
  --nios2_fpu_burst_5_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_5_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_5_upstream_begins_xfer) = '1' then 
        nios2_fpu_burst_5_upstream_reg_firsttransfer <= nios2_fpu_burst_5_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_5_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  nios2_fpu_burst_5_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_nios2_fpu_burst_5_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_5_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_nios2_fpu_burst_5_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_nios2_fpu_burst_5_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_5_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (nios2_fpu_burst_5_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --nios2_fpu_burst_5_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_5_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_5_upstream_begins_xfer) = '1' then 
        nios2_fpu_burst_5_upstream_bbt_burstcounter <= nios2_fpu_burst_5_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_5_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_fpu_burst_5_upstream_beginbursttransfer_internal <= nios2_fpu_burst_5_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_5_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --nios2_fpu_burst_5_upstream_read assignment, which is an e_mux
  internal_nios2_fpu_burst_5_upstream_read <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream AND nios2_fast_fpu_data_master_read;
  --nios2_fpu_burst_5_upstream_write assignment, which is an e_mux
  internal_nios2_fpu_burst_5_upstream_write <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream AND nios2_fast_fpu_data_master_write;
  --nios2_fpu_burst_5_upstream_address mux, which is an e_mux
  nios2_fpu_burst_5_upstream_address <= nios2_fast_fpu_data_master_address_to_slave (10 DOWNTO 0);
  --d1_nios2_fpu_burst_5_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_fpu_burst_5_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_fpu_burst_5_upstream_end_xfer <= nios2_fpu_burst_5_upstream_end_xfer;
    end if;

  end process;

  --nios2_fpu_burst_5_upstream_waits_for_read in a cycle, which is an e_mux
  nios2_fpu_burst_5_upstream_waits_for_read <= nios2_fpu_burst_5_upstream_in_a_read_cycle AND internal_nios2_fpu_burst_5_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_5_upstream_in_a_read_cycle assignment, which is an e_assign
  nios2_fpu_burst_5_upstream_in_a_read_cycle <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream AND nios2_fast_fpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_fpu_burst_5_upstream_in_a_read_cycle;
  --nios2_fpu_burst_5_upstream_waits_for_write in a cycle, which is an e_mux
  nios2_fpu_burst_5_upstream_waits_for_write <= nios2_fpu_burst_5_upstream_in_a_write_cycle AND internal_nios2_fpu_burst_5_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_5_upstream_in_a_write_cycle assignment, which is an e_assign
  nios2_fpu_burst_5_upstream_in_a_write_cycle <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream AND nios2_fast_fpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_fpu_burst_5_upstream_in_a_write_cycle;
  wait_for_nios2_fpu_burst_5_upstream_counter <= std_logic'('0');
  --nios2_fpu_burst_5_upstream_byteenable byte enable port mux, which is an e_mux
  nios2_fpu_burst_5_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --burstcount mux, which is an e_mux
  internal_nios2_fpu_burst_5_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  nios2_fpu_burst_5_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream;
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream <= internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream;
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream <= internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream;
  --vhdl renameroo for output signals
  nios2_fpu_burst_5_upstream_burstcount <= internal_nios2_fpu_burst_5_upstream_burstcount;
  --vhdl renameroo for output signals
  nios2_fpu_burst_5_upstream_read <= internal_nios2_fpu_burst_5_upstream_read;
  --vhdl renameroo for output signals
  nios2_fpu_burst_5_upstream_waitrequest_from_sa <= internal_nios2_fpu_burst_5_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  nios2_fpu_burst_5_upstream_write <= internal_nios2_fpu_burst_5_upstream_write;
--synthesis translate_off
    --nios2_fpu_burst_5/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --nios2_fast_fpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line61 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line61, now);
          write(write_line61, string'(": "));
          write(write_line61, string'("nios2_fast_fpu/data_master drove 0 on its 'burstcount' port while accessing slave nios2_fpu_burst_5/upstream"));
          write(output, write_line61.all);
          deallocate (write_line61);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_5_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_nios2_fast_fpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal nios2_fast_fpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_5_downstream_address : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal nios2_fpu_burst_5_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_fpu_burst_5_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal nios2_fpu_burst_5_downstream_latency_counter : OUT STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_5_downstream_readdatavalid : OUT STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_reset_n : OUT STD_LOGIC;
                 signal nios2_fpu_burst_5_downstream_waitrequest : OUT STD_LOGIC
              );
end entity nios2_fpu_burst_5_downstream_arbitrator;


architecture europa of nios2_fpu_burst_5_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_fpu_burst_5_downstream_address_to_slave :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal internal_nios2_fpu_burst_5_downstream_latency_counter :  STD_LOGIC;
                signal internal_nios2_fpu_burst_5_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_address_last_time :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_5_downstream_burstcount_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_5_downstream_is_granted_some_slave :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_read_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_run :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_write_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_nios2_fpu_burst_5_downstream_latency_counter :  STD_LOGIC;
                signal pre_flush_nios2_fpu_burst_5_downstream_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module OR NOT nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module OR NOT nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module OR NOT nios2_fpu_burst_5_downstream_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_nios2_fast_fpu_jtag_debug_module_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_5_downstream_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module OR NOT nios2_fpu_burst_5_downstream_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_5_downstream_write)))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_fpu_burst_5_downstream_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_fpu_burst_5_downstream_address_to_slave <= nios2_fpu_burst_5_downstream_address;
  --nios2_fpu_burst_5_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_5_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      nios2_fpu_burst_5_downstream_read_but_no_slave_selected <= (nios2_fpu_burst_5_downstream_read AND nios2_fpu_burst_5_downstream_run) AND NOT nios2_fpu_burst_5_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  nios2_fpu_burst_5_downstream_is_granted_some_slave <= nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_nios2_fpu_burst_5_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  nios2_fpu_burst_5_downstream_readdatavalid <= (nios2_fpu_burst_5_downstream_read_but_no_slave_selected OR pre_flush_nios2_fpu_burst_5_downstream_readdatavalid) OR nios2_fpu_burst_5_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module;
  --nios2_fpu_burst_5/downstream readdata mux, which is an e_mux
  nios2_fpu_burst_5_downstream_readdata <= nios2_fast_fpu_jtag_debug_module_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_fpu_burst_5_downstream_waitrequest <= NOT nios2_fpu_burst_5_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_nios2_fpu_burst_5_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_nios2_fpu_burst_5_downstream_latency_counter <= p1_nios2_fpu_burst_5_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_nios2_fpu_burst_5_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((nios2_fpu_burst_5_downstream_run AND nios2_fpu_burst_5_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_5_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_5_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --nios2_fpu_burst_5_downstream_reset_n assignment, which is an e_assign
  nios2_fpu_burst_5_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_fpu_burst_5_downstream_address_to_slave <= internal_nios2_fpu_burst_5_downstream_address_to_slave;
  --vhdl renameroo for output signals
  nios2_fpu_burst_5_downstream_latency_counter <= internal_nios2_fpu_burst_5_downstream_latency_counter;
  --vhdl renameroo for output signals
  nios2_fpu_burst_5_downstream_waitrequest <= internal_nios2_fpu_burst_5_downstream_waitrequest;
--synthesis translate_off
    --nios2_fpu_burst_5_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_5_downstream_address_last_time <= std_logic_vector'("00000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_5_downstream_address_last_time <= nios2_fpu_burst_5_downstream_address;
      end if;

    end process;

    --nios2_fpu_burst_5/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_fpu_burst_5_downstream_waitrequest AND ((nios2_fpu_burst_5_downstream_read OR nios2_fpu_burst_5_downstream_write));
      end if;

    end process;

    --nios2_fpu_burst_5_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line62 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_5_downstream_address /= nios2_fpu_burst_5_downstream_address_last_time))))) = '1' then 
          write(write_line62, now);
          write(write_line62, string'(": "));
          write(write_line62, string'("nios2_fpu_burst_5_downstream_address did not heed wait!!!"));
          write(output, write_line62.all);
          deallocate (write_line62);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_5_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_5_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_5_downstream_burstcount_last_time <= nios2_fpu_burst_5_downstream_burstcount;
      end if;

    end process;

    --nios2_fpu_burst_5_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line63 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_5_downstream_burstcount) /= std_logic'(nios2_fpu_burst_5_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line63, now);
          write(write_line63, string'(": "));
          write(write_line63, string'("nios2_fpu_burst_5_downstream_burstcount did not heed wait!!!"));
          write(output, write_line63.all);
          deallocate (write_line63);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_5_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_5_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_5_downstream_byteenable_last_time <= nios2_fpu_burst_5_downstream_byteenable;
      end if;

    end process;

    --nios2_fpu_burst_5_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line64 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_5_downstream_byteenable /= nios2_fpu_burst_5_downstream_byteenable_last_time))))) = '1' then 
          write(write_line64, now);
          write(write_line64, string'(": "));
          write(write_line64, string'("nios2_fpu_burst_5_downstream_byteenable did not heed wait!!!"));
          write(output, write_line64.all);
          deallocate (write_line64);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_5_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_5_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_5_downstream_read_last_time <= nios2_fpu_burst_5_downstream_read;
      end if;

    end process;

    --nios2_fpu_burst_5_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line65 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_5_downstream_read) /= std_logic'(nios2_fpu_burst_5_downstream_read_last_time)))))) = '1' then 
          write(write_line65, now);
          write(write_line65, string'(": "));
          write(write_line65, string'("nios2_fpu_burst_5_downstream_read did not heed wait!!!"));
          write(output, write_line65.all);
          deallocate (write_line65);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_5_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_5_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_5_downstream_write_last_time <= nios2_fpu_burst_5_downstream_write;
      end if;

    end process;

    --nios2_fpu_burst_5_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line66 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_5_downstream_write) /= std_logic'(nios2_fpu_burst_5_downstream_write_last_time)))))) = '1' then 
          write(write_line66, now);
          write(write_line66, string'(": "));
          write(write_line66, string'("nios2_fpu_burst_5_downstream_write did not heed wait!!!"));
          write(output, write_line66.all);
          deallocate (write_line66);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_5_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_5_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_5_downstream_writedata_last_time <= nios2_fpu_burst_5_downstream_writedata;
      end if;

    end process;

    --nios2_fpu_burst_5_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line67 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_5_downstream_writedata /= nios2_fpu_burst_5_downstream_writedata_last_time)))) AND nios2_fpu_burst_5_downstream_write)) = '1' then 
          write(write_line67, now);
          write(write_line67, string'(": "));
          write(write_line67, string'("nios2_fpu_burst_5_downstream_writedata did not heed wait!!!"));
          write(output, write_line67.all);
          deallocate (write_line67);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_nios2_fpu_burst_6_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_nios2_fpu_burst_6_upstream_module;


architecture europa of burstcount_fifo_for_nios2_fpu_burst_6_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_2;
  empty <= NOT(full_0);
  full_3 <= std_logic'('0');
  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("0000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_6_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_6_upstream_module;


architecture europa of rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_6_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_2;
  empty <= NOT(full_0);
  full_3 <= std_logic'('0');
  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_6_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_debugaccess : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_latency_counter : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_write : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_6_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_6_upstream_readdatavalid : IN STD_LOGIC;
                 signal nios2_fpu_burst_6_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_nios2_fpu_burst_6_upstream_end_xfer : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream : OUT STD_LOGIC;
                 signal nios2_fpu_burst_6_upstream_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_burst_6_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_6_upstream_byteaddress : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                 signal nios2_fpu_burst_6_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_6_upstream_debugaccess : OUT STD_LOGIC;
                 signal nios2_fpu_burst_6_upstream_read : OUT STD_LOGIC;
                 signal nios2_fpu_burst_6_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_6_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_fpu_burst_6_upstream_write : OUT STD_LOGIC;
                 signal nios2_fpu_burst_6_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity nios2_fpu_burst_6_upstream_arbitrator;


architecture europa of nios2_fpu_burst_6_upstream_arbitrator is
component burstcount_fifo_for_nios2_fpu_burst_6_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_nios2_fpu_burst_6_upstream_module;

component rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_6_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_6_upstream_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_fpu_burst_6_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream :  STD_LOGIC;
                signal internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream :  STD_LOGIC;
                signal internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream :  STD_LOGIC;
                signal internal_nios2_fpu_burst_6_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_nios2_fpu_burst_6_upstream_read :  STD_LOGIC;
                signal internal_nios2_fpu_burst_6_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_nios2_fpu_burst_6_upstream_write :  STD_LOGIC;
                signal module_input36 :  STD_LOGIC;
                signal module_input37 :  STD_LOGIC;
                signal module_input38 :  STD_LOGIC;
                signal module_input39 :  STD_LOGIC;
                signal module_input40 :  STD_LOGIC;
                signal module_input41 :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_arbiterlock :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_continuerequest :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_rdv_fifo_empty_nios2_fpu_burst_6_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_rdv_fifo_output_from_nios2_fpu_burst_6_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_saved_grant_nios2_fpu_burst_6_upstream :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_allgrants :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_any_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_arb_counter_enable :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_arb_share_counter :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_begins_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_end_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_grant_vector :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_in_a_read_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_in_a_write_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_load_fifo :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_master_qreq_vector :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_reg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_waits_for_read :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_waits_for_write :  STD_LOGIC;
                signal p0_nios2_fpu_burst_6_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_nios2_fpu_burst_6_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_fpu_burst_6_upstream_end_xfer;
    end if;

  end process;

  nios2_fpu_burst_6_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream);
  --assign nios2_fpu_burst_6_upstream_readdatavalid_from_sa = nios2_fpu_burst_6_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_6_upstream_readdatavalid_from_sa <= nios2_fpu_burst_6_upstream_readdatavalid;
  --assign nios2_fpu_burst_6_upstream_readdata_from_sa = nios2_fpu_burst_6_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_6_upstream_readdata_from_sa <= nios2_fpu_burst_6_upstream_readdata;
  internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream <= to_std_logic(((Std_Logic_Vector'(nios2_fast_fpu_data_master_address_to_slave(28 DOWNTO 13) & std_logic_vector'("0000000000000")) = std_logic_vector'("01111000000000000000000000000")))) AND ((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write));
  --assign nios2_fpu_burst_6_upstream_waitrequest_from_sa = nios2_fpu_burst_6_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_fpu_burst_6_upstream_waitrequest_from_sa <= nios2_fpu_burst_6_upstream_waitrequest;
  --nios2_fpu_burst_6_upstream_arb_share_counter set values, which is an e_mux
  nios2_fpu_burst_6_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((nios2_fast_fpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 6);
  --nios2_fpu_burst_6_upstream_non_bursting_master_requests mux, which is an e_mux
  nios2_fpu_burst_6_upstream_non_bursting_master_requests <= std_logic'('0');
  --nios2_fpu_burst_6_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_fpu_burst_6_upstream_any_bursting_master_saved_grant <= nios2_fast_fpu_data_master_saved_grant_nios2_fpu_burst_6_upstream;
  --nios2_fpu_burst_6_upstream_arb_share_counter_next_value assignment, which is an e_assign
  nios2_fpu_burst_6_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_6_upstream_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_6_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_fpu_burst_6_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_6_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 6);
  --nios2_fpu_burst_6_upstream_allgrants all slave grants, which is an e_mux
  nios2_fpu_burst_6_upstream_allgrants <= nios2_fpu_burst_6_upstream_grant_vector;
  --nios2_fpu_burst_6_upstream_end_xfer assignment, which is an e_assign
  nios2_fpu_burst_6_upstream_end_xfer <= NOT ((nios2_fpu_burst_6_upstream_waits_for_read OR nios2_fpu_burst_6_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_fpu_burst_6_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_fpu_burst_6_upstream <= nios2_fpu_burst_6_upstream_end_xfer AND (((NOT nios2_fpu_burst_6_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_fpu_burst_6_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_fpu_burst_6_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_fpu_burst_6_upstream AND nios2_fpu_burst_6_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_6_upstream AND NOT nios2_fpu_burst_6_upstream_non_bursting_master_requests));
  --nios2_fpu_burst_6_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_6_upstream_arb_share_counter <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_6_upstream_arb_counter_enable) = '1' then 
        nios2_fpu_burst_6_upstream_arb_share_counter <= nios2_fpu_burst_6_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_6_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_6_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_fpu_burst_6_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_fpu_burst_6_upstream)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_6_upstream AND NOT nios2_fpu_burst_6_upstream_non_bursting_master_requests)))) = '1' then 
        nios2_fpu_burst_6_upstream_slavearbiterlockenable <= or_reduce(nios2_fpu_burst_6_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --nios2_fast_fpu/data_master nios2_fpu_burst_6/upstream arbiterlock, which is an e_assign
  nios2_fast_fpu_data_master_arbiterlock <= nios2_fpu_burst_6_upstream_slavearbiterlockenable AND nios2_fast_fpu_data_master_continuerequest;
  --nios2_fpu_burst_6_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_fpu_burst_6_upstream_slavearbiterlockenable2 <= or_reduce(nios2_fpu_burst_6_upstream_arb_share_counter_next_value);
  --nios2_fast_fpu/data_master nios2_fpu_burst_6/upstream arbiterlock2, which is an e_assign
  nios2_fast_fpu_data_master_arbiterlock2 <= nios2_fpu_burst_6_upstream_slavearbiterlockenable2 AND nios2_fast_fpu_data_master_continuerequest;
  --nios2_fpu_burst_6_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_fpu_burst_6_upstream_any_continuerequest <= std_logic'('1');
  --nios2_fast_fpu_data_master_continuerequest continued request, which is an e_assign
  nios2_fast_fpu_data_master_continuerequest <= std_logic'('1');
  internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream <= internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream AND NOT ((nios2_fast_fpu_data_master_read AND ((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_data_master_latency_counter))))))) OR (nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register)) OR (nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register)) OR (nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register)))));
  --unique name for nios2_fpu_burst_6_upstream_move_on_to_next_transaction, which is an e_assign
  nios2_fpu_burst_6_upstream_move_on_to_next_transaction <= nios2_fpu_burst_6_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_6_upstream_load_fifo;
  --the currently selected burstcount for nios2_fpu_burst_6_upstream, which is an e_mux
  nios2_fpu_burst_6_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_nios2_fpu_burst_6_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_nios2_fpu_burst_6_upstream : burstcount_fifo_for_nios2_fpu_burst_6_upstream_module
    port map(
      data_out => nios2_fpu_burst_6_upstream_transaction_burst_count,
      empty => nios2_fpu_burst_6_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input36,
      clk => clk,
      data_in => nios2_fpu_burst_6_upstream_selected_burstcount,
      read => nios2_fpu_burst_6_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input37,
      write => module_input38
    );

  module_input36 <= std_logic'('0');
  module_input37 <= std_logic'('0');
  module_input38 <= ((in_a_read_cycle AND NOT nios2_fpu_burst_6_upstream_waits_for_read) AND nios2_fpu_burst_6_upstream_load_fifo) AND NOT ((nios2_fpu_burst_6_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_6_upstream_burstcount_fifo_empty));

  --nios2_fpu_burst_6_upstream current burst minus one, which is an e_assign
  nios2_fpu_burst_6_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_6_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for nios2_fpu_burst_6_upstream, which is an e_mux
  nios2_fpu_burst_6_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_6_upstream_waits_for_read)) AND NOT nios2_fpu_burst_6_upstream_load_fifo))) = '1'), nios2_fpu_burst_6_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_6_upstream_waits_for_read) AND nios2_fpu_burst_6_upstream_this_cycle_is_the_last_burst) AND nios2_fpu_burst_6_upstream_burstcount_fifo_empty))) = '1'), nios2_fpu_burst_6_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((nios2_fpu_burst_6_upstream_this_cycle_is_the_last_burst)) = '1'), nios2_fpu_burst_6_upstream_transaction_burst_count, nios2_fpu_burst_6_upstream_current_burst_minus_one)));
  --the current burst count for nios2_fpu_burst_6_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_6_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((nios2_fpu_burst_6_upstream_readdatavalid_from_sa OR ((NOT nios2_fpu_burst_6_upstream_load_fifo AND ((in_a_read_cycle AND NOT nios2_fpu_burst_6_upstream_waits_for_read)))))) = '1' then 
        nios2_fpu_burst_6_upstream_current_burst <= nios2_fpu_burst_6_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_nios2_fpu_burst_6_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT nios2_fpu_burst_6_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_6_upstream_waits_for_read)) AND nios2_fpu_burst_6_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_6_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_6_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_6_upstream_waits_for_read)) AND NOT nios2_fpu_burst_6_upstream_load_fifo) OR nios2_fpu_burst_6_upstream_this_cycle_is_the_last_burst)) = '1' then 
        nios2_fpu_burst_6_upstream_load_fifo <= p0_nios2_fpu_burst_6_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for nios2_fpu_burst_6_upstream, which is an e_assign
  nios2_fpu_burst_6_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(nios2_fpu_burst_6_upstream_current_burst_minus_one)) AND nios2_fpu_burst_6_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_6_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_6_upstream : rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_6_upstream_module
    port map(
      data_out => nios2_fast_fpu_data_master_rdv_fifo_output_from_nios2_fpu_burst_6_upstream,
      empty => open,
      fifo_contains_ones_n => nios2_fast_fpu_data_master_rdv_fifo_empty_nios2_fpu_burst_6_upstream,
      full => open,
      clear_fifo => module_input39,
      clk => clk,
      data_in => internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream,
      read => nios2_fpu_burst_6_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input40,
      write => module_input41
    );

  module_input39 <= std_logic'('0');
  module_input40 <= std_logic'('0');
  module_input41 <= in_a_read_cycle AND NOT nios2_fpu_burst_6_upstream_waits_for_read;

  nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register <= NOT nios2_fast_fpu_data_master_rdv_fifo_empty_nios2_fpu_burst_6_upstream;
  --local readdatavalid nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream, which is an e_mux
  nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream <= nios2_fpu_burst_6_upstream_readdatavalid_from_sa;
  --nios2_fpu_burst_6_upstream_writedata mux, which is an e_mux
  nios2_fpu_burst_6_upstream_writedata <= nios2_fast_fpu_data_master_writedata;
  --byteaddress mux for nios2_fpu_burst_6/upstream, which is an e_mux
  nios2_fpu_burst_6_upstream_byteaddress <= nios2_fast_fpu_data_master_address_to_slave (14 DOWNTO 0);
  --master is always granted when requested
  internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream <= internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream;
  --nios2_fast_fpu/data_master saved-grant nios2_fpu_burst_6/upstream, which is an e_assign
  nios2_fast_fpu_data_master_saved_grant_nios2_fpu_burst_6_upstream <= internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream;
  --allow new arb cycle for nios2_fpu_burst_6/upstream, which is an e_assign
  nios2_fpu_burst_6_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_fpu_burst_6_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_fpu_burst_6_upstream_master_qreq_vector <= std_logic'('1');
  --nios2_fpu_burst_6_upstream_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_6_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_fpu_burst_6_upstream_begins_xfer) = '1'), nios2_fpu_burst_6_upstream_unreg_firsttransfer, nios2_fpu_burst_6_upstream_reg_firsttransfer);
  --nios2_fpu_burst_6_upstream_unreg_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_6_upstream_unreg_firsttransfer <= NOT ((nios2_fpu_burst_6_upstream_slavearbiterlockenable AND nios2_fpu_burst_6_upstream_any_continuerequest));
  --nios2_fpu_burst_6_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_6_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_6_upstream_begins_xfer) = '1' then 
        nios2_fpu_burst_6_upstream_reg_firsttransfer <= nios2_fpu_burst_6_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_6_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  nios2_fpu_burst_6_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_nios2_fpu_burst_6_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_6_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_nios2_fpu_burst_6_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_nios2_fpu_burst_6_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_6_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (nios2_fpu_burst_6_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --nios2_fpu_burst_6_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_6_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_6_upstream_begins_xfer) = '1' then 
        nios2_fpu_burst_6_upstream_bbt_burstcounter <= nios2_fpu_burst_6_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_6_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_fpu_burst_6_upstream_beginbursttransfer_internal <= nios2_fpu_burst_6_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_6_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --nios2_fpu_burst_6_upstream_read assignment, which is an e_mux
  internal_nios2_fpu_burst_6_upstream_read <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream AND nios2_fast_fpu_data_master_read;
  --nios2_fpu_burst_6_upstream_write assignment, which is an e_mux
  internal_nios2_fpu_burst_6_upstream_write <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream AND nios2_fast_fpu_data_master_write;
  --nios2_fpu_burst_6_upstream_address mux, which is an e_mux
  nios2_fpu_burst_6_upstream_address <= nios2_fast_fpu_data_master_address_to_slave (12 DOWNTO 0);
  --d1_nios2_fpu_burst_6_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_fpu_burst_6_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_fpu_burst_6_upstream_end_xfer <= nios2_fpu_burst_6_upstream_end_xfer;
    end if;

  end process;

  --nios2_fpu_burst_6_upstream_waits_for_read in a cycle, which is an e_mux
  nios2_fpu_burst_6_upstream_waits_for_read <= nios2_fpu_burst_6_upstream_in_a_read_cycle AND internal_nios2_fpu_burst_6_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_6_upstream_in_a_read_cycle assignment, which is an e_assign
  nios2_fpu_burst_6_upstream_in_a_read_cycle <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream AND nios2_fast_fpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_fpu_burst_6_upstream_in_a_read_cycle;
  --nios2_fpu_burst_6_upstream_waits_for_write in a cycle, which is an e_mux
  nios2_fpu_burst_6_upstream_waits_for_write <= nios2_fpu_burst_6_upstream_in_a_write_cycle AND internal_nios2_fpu_burst_6_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_6_upstream_in_a_write_cycle assignment, which is an e_assign
  nios2_fpu_burst_6_upstream_in_a_write_cycle <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream AND nios2_fast_fpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_fpu_burst_6_upstream_in_a_write_cycle;
  wait_for_nios2_fpu_burst_6_upstream_counter <= std_logic'('0');
  --nios2_fpu_burst_6_upstream_byteenable byte enable port mux, which is an e_mux
  nios2_fpu_burst_6_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --burstcount mux, which is an e_mux
  internal_nios2_fpu_burst_6_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  nios2_fpu_burst_6_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream;
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream <= internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream;
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream <= internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream;
  --vhdl renameroo for output signals
  nios2_fpu_burst_6_upstream_burstcount <= internal_nios2_fpu_burst_6_upstream_burstcount;
  --vhdl renameroo for output signals
  nios2_fpu_burst_6_upstream_read <= internal_nios2_fpu_burst_6_upstream_read;
  --vhdl renameroo for output signals
  nios2_fpu_burst_6_upstream_waitrequest_from_sa <= internal_nios2_fpu_burst_6_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  nios2_fpu_burst_6_upstream_write <= internal_nios2_fpu_burst_6_upstream_write;
--synthesis translate_off
    --nios2_fpu_burst_6/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --nios2_fast_fpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line68 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line68, now);
          write(write_line68, string'(": "));
          write(write_line68, string'("nios2_fast_fpu/data_master drove 0 on its 'burstcount' port while accessing slave nios2_fpu_burst_6/upstream"));
          write(output, write_line68.all);
          deallocate (write_line68);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_6_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_ipl_memory_s1_end_xfer : IN STD_LOGIC;
                 signal ipl_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_6_downstream_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_burst_6_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_requests_ipl_memory_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_fpu_burst_6_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_burst_6_downstream_latency_counter : OUT STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_6_downstream_readdatavalid : OUT STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_reset_n : OUT STD_LOGIC;
                 signal nios2_fpu_burst_6_downstream_waitrequest : OUT STD_LOGIC
              );
end entity nios2_fpu_burst_6_downstream_arbitrator;


architecture europa of nios2_fpu_burst_6_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_fpu_burst_6_downstream_address_to_slave :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal internal_nios2_fpu_burst_6_downstream_latency_counter :  STD_LOGIC;
                signal internal_nios2_fpu_burst_6_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_address_last_time :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_6_downstream_burstcount_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_6_downstream_is_granted_some_slave :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_read_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_run :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_write_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_nios2_fpu_burst_6_downstream_latency_counter :  STD_LOGIC;
                signal pre_flush_nios2_fpu_burst_6_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1 OR NOT nios2_fpu_burst_6_downstream_requests_ipl_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 OR NOT nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1 OR NOT ((nios2_fpu_burst_6_downstream_read OR nios2_fpu_burst_6_downstream_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_6_downstream_read OR nios2_fpu_burst_6_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1 OR NOT ((nios2_fpu_burst_6_downstream_read OR nios2_fpu_burst_6_downstream_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_6_downstream_read OR nios2_fpu_burst_6_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_fpu_burst_6_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_fpu_burst_6_downstream_address_to_slave <= nios2_fpu_burst_6_downstream_address;
  --nios2_fpu_burst_6_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_6_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      nios2_fpu_burst_6_downstream_read_but_no_slave_selected <= (nios2_fpu_burst_6_downstream_read AND nios2_fpu_burst_6_downstream_run) AND NOT nios2_fpu_burst_6_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  nios2_fpu_burst_6_downstream_is_granted_some_slave <= nios2_fpu_burst_6_downstream_granted_ipl_memory_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_nios2_fpu_burst_6_downstream_readdatavalid <= nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  nios2_fpu_burst_6_downstream_readdatavalid <= nios2_fpu_burst_6_downstream_read_but_no_slave_selected OR pre_flush_nios2_fpu_burst_6_downstream_readdatavalid;
  --nios2_fpu_burst_6/downstream readdata mux, which is an e_mux
  nios2_fpu_burst_6_downstream_readdata <= ipl_memory_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_fpu_burst_6_downstream_waitrequest <= NOT nios2_fpu_burst_6_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_nios2_fpu_burst_6_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_nios2_fpu_burst_6_downstream_latency_counter <= p1_nios2_fpu_burst_6_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_nios2_fpu_burst_6_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((nios2_fpu_burst_6_downstream_run AND nios2_fpu_burst_6_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_6_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_6_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_6_downstream_requests_ipl_memory_s1))) AND std_logic_vector'("00000000000000000000000000000001")));
  --nios2_fpu_burst_6_downstream_reset_n assignment, which is an e_assign
  nios2_fpu_burst_6_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_fpu_burst_6_downstream_address_to_slave <= internal_nios2_fpu_burst_6_downstream_address_to_slave;
  --vhdl renameroo for output signals
  nios2_fpu_burst_6_downstream_latency_counter <= internal_nios2_fpu_burst_6_downstream_latency_counter;
  --vhdl renameroo for output signals
  nios2_fpu_burst_6_downstream_waitrequest <= internal_nios2_fpu_burst_6_downstream_waitrequest;
--synthesis translate_off
    --nios2_fpu_burst_6_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_6_downstream_address_last_time <= std_logic_vector'("0000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_6_downstream_address_last_time <= nios2_fpu_burst_6_downstream_address;
      end if;

    end process;

    --nios2_fpu_burst_6/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_fpu_burst_6_downstream_waitrequest AND ((nios2_fpu_burst_6_downstream_read OR nios2_fpu_burst_6_downstream_write));
      end if;

    end process;

    --nios2_fpu_burst_6_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line69 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_6_downstream_address /= nios2_fpu_burst_6_downstream_address_last_time))))) = '1' then 
          write(write_line69, now);
          write(write_line69, string'(": "));
          write(write_line69, string'("nios2_fpu_burst_6_downstream_address did not heed wait!!!"));
          write(output, write_line69.all);
          deallocate (write_line69);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_6_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_6_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_6_downstream_burstcount_last_time <= nios2_fpu_burst_6_downstream_burstcount;
      end if;

    end process;

    --nios2_fpu_burst_6_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line70 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_6_downstream_burstcount) /= std_logic'(nios2_fpu_burst_6_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line70, now);
          write(write_line70, string'(": "));
          write(write_line70, string'("nios2_fpu_burst_6_downstream_burstcount did not heed wait!!!"));
          write(output, write_line70.all);
          deallocate (write_line70);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_6_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_6_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_6_downstream_byteenable_last_time <= nios2_fpu_burst_6_downstream_byteenable;
      end if;

    end process;

    --nios2_fpu_burst_6_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line71 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_6_downstream_byteenable /= nios2_fpu_burst_6_downstream_byteenable_last_time))))) = '1' then 
          write(write_line71, now);
          write(write_line71, string'(": "));
          write(write_line71, string'("nios2_fpu_burst_6_downstream_byteenable did not heed wait!!!"));
          write(output, write_line71.all);
          deallocate (write_line71);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_6_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_6_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_6_downstream_read_last_time <= nios2_fpu_burst_6_downstream_read;
      end if;

    end process;

    --nios2_fpu_burst_6_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line72 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_6_downstream_read) /= std_logic'(nios2_fpu_burst_6_downstream_read_last_time)))))) = '1' then 
          write(write_line72, now);
          write(write_line72, string'(": "));
          write(write_line72, string'("nios2_fpu_burst_6_downstream_read did not heed wait!!!"));
          write(output, write_line72.all);
          deallocate (write_line72);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_6_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_6_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_6_downstream_write_last_time <= nios2_fpu_burst_6_downstream_write;
      end if;

    end process;

    --nios2_fpu_burst_6_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line73 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_6_downstream_write) /= std_logic'(nios2_fpu_burst_6_downstream_write_last_time)))))) = '1' then 
          write(write_line73, now);
          write(write_line73, string'(": "));
          write(write_line73, string'("nios2_fpu_burst_6_downstream_write did not heed wait!!!"));
          write(output, write_line73.all);
          deallocate (write_line73);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_6_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_6_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_6_downstream_writedata_last_time <= nios2_fpu_burst_6_downstream_writedata;
      end if;

    end process;

    --nios2_fpu_burst_6_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line74 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_6_downstream_writedata /= nios2_fpu_burst_6_downstream_writedata_last_time)))) AND nios2_fpu_burst_6_downstream_write)) = '1' then 
          write(write_line74, now);
          write(write_line74, string'(": "));
          write(write_line74, string'("nios2_fpu_burst_6_downstream_writedata did not heed wait!!!"));
          write(output, write_line74.all);
          deallocate (write_line74);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_nios2_fpu_burst_7_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_nios2_fpu_burst_7_upstream_module;


architecture europa of burstcount_fifo_for_nios2_fpu_burst_7_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_2;
  empty <= NOT(full_0);
  full_3 <= std_logic'('0');
  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("0000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_7_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_7_upstream_module;


architecture europa of rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_7_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_2;
  empty <= NOT(full_0);
  full_3 <= std_logic'('0');
  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_7_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal nios2_fast_fpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fast_fpu_instruction_master_latency_counter : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fpu_burst_7_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_7_upstream_readdatavalid : IN STD_LOGIC;
                 signal nios2_fpu_burst_7_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_nios2_fpu_burst_7_upstream_end_xfer : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register : OUT STD_LOGIC;
                 signal nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream : OUT STD_LOGIC;
                 signal nios2_fpu_burst_7_upstream_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_burst_7_upstream_byteaddress : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                 signal nios2_fpu_burst_7_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_7_upstream_debugaccess : OUT STD_LOGIC;
                 signal nios2_fpu_burst_7_upstream_read : OUT STD_LOGIC;
                 signal nios2_fpu_burst_7_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_7_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_fpu_burst_7_upstream_write : OUT STD_LOGIC
              );
end entity nios2_fpu_burst_7_upstream_arbitrator;


architecture europa of nios2_fpu_burst_7_upstream_arbitrator is
component burstcount_fifo_for_nios2_fpu_burst_7_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_nios2_fpu_burst_7_upstream_module;

component rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_7_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_7_upstream_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_fpu_burst_7_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream :  STD_LOGIC;
                signal internal_nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream :  STD_LOGIC;
                signal internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream :  STD_LOGIC;
                signal internal_nios2_fpu_burst_7_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal module_input42 :  STD_LOGIC;
                signal module_input43 :  STD_LOGIC;
                signal module_input44 :  STD_LOGIC;
                signal module_input45 :  STD_LOGIC;
                signal module_input46 :  STD_LOGIC;
                signal module_input47 :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_continuerequest :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_rdv_fifo_empty_nios2_fpu_burst_7_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_rdv_fifo_output_from_nios2_fpu_burst_7_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_saved_grant_nios2_fpu_burst_7_upstream :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_allgrants :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_any_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_arb_counter_enable :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_arb_share_counter :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_7_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_7_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_7_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_begins_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_7_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_7_upstream_end_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_grant_vector :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_in_a_read_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_in_a_write_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_load_fifo :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_master_qreq_vector :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_7_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_reg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_7_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_7_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_waits_for_read :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_waits_for_write :  STD_LOGIC;
                signal p0_nios2_fpu_burst_7_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_nios2_fpu_burst_7_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_fpu_burst_7_upstream_end_xfer;
    end if;

  end process;

  nios2_fpu_burst_7_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream);
  --assign nios2_fpu_burst_7_upstream_readdatavalid_from_sa = nios2_fpu_burst_7_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_7_upstream_readdatavalid_from_sa <= nios2_fpu_burst_7_upstream_readdatavalid;
  --assign nios2_fpu_burst_7_upstream_readdata_from_sa = nios2_fpu_burst_7_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_7_upstream_readdata_from_sa <= nios2_fpu_burst_7_upstream_readdata;
  internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream <= ((to_std_logic(((Std_Logic_Vector'(nios2_fast_fpu_instruction_master_address_to_slave(27 DOWNTO 13) & std_logic_vector'("0000000000000")) = std_logic_vector'("1111000000000000000000000000")))) AND (nios2_fast_fpu_instruction_master_read))) AND nios2_fast_fpu_instruction_master_read;
  --assign nios2_fpu_burst_7_upstream_waitrequest_from_sa = nios2_fpu_burst_7_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_fpu_burst_7_upstream_waitrequest_from_sa <= nios2_fpu_burst_7_upstream_waitrequest;
  --nios2_fpu_burst_7_upstream_arb_share_counter set values, which is an e_mux
  nios2_fpu_burst_7_upstream_arb_share_set_values <= std_logic_vector'("000001");
  --nios2_fpu_burst_7_upstream_non_bursting_master_requests mux, which is an e_mux
  nios2_fpu_burst_7_upstream_non_bursting_master_requests <= std_logic'('0');
  --nios2_fpu_burst_7_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_fpu_burst_7_upstream_any_bursting_master_saved_grant <= nios2_fast_fpu_instruction_master_saved_grant_nios2_fpu_burst_7_upstream;
  --nios2_fpu_burst_7_upstream_arb_share_counter_next_value assignment, which is an e_assign
  nios2_fpu_burst_7_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_7_upstream_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_7_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_fpu_burst_7_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_7_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 6);
  --nios2_fpu_burst_7_upstream_allgrants all slave grants, which is an e_mux
  nios2_fpu_burst_7_upstream_allgrants <= nios2_fpu_burst_7_upstream_grant_vector;
  --nios2_fpu_burst_7_upstream_end_xfer assignment, which is an e_assign
  nios2_fpu_burst_7_upstream_end_xfer <= NOT ((nios2_fpu_burst_7_upstream_waits_for_read OR nios2_fpu_burst_7_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_fpu_burst_7_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_fpu_burst_7_upstream <= nios2_fpu_burst_7_upstream_end_xfer AND (((NOT nios2_fpu_burst_7_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_fpu_burst_7_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_fpu_burst_7_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_fpu_burst_7_upstream AND nios2_fpu_burst_7_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_7_upstream AND NOT nios2_fpu_burst_7_upstream_non_bursting_master_requests));
  --nios2_fpu_burst_7_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_7_upstream_arb_share_counter <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_7_upstream_arb_counter_enable) = '1' then 
        nios2_fpu_burst_7_upstream_arb_share_counter <= nios2_fpu_burst_7_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_7_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_7_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_fpu_burst_7_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_fpu_burst_7_upstream)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_7_upstream AND NOT nios2_fpu_burst_7_upstream_non_bursting_master_requests)))) = '1' then 
        nios2_fpu_burst_7_upstream_slavearbiterlockenable <= or_reduce(nios2_fpu_burst_7_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --nios2_fast_fpu/instruction_master nios2_fpu_burst_7/upstream arbiterlock, which is an e_assign
  nios2_fast_fpu_instruction_master_arbiterlock <= nios2_fpu_burst_7_upstream_slavearbiterlockenable AND nios2_fast_fpu_instruction_master_continuerequest;
  --nios2_fpu_burst_7_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_fpu_burst_7_upstream_slavearbiterlockenable2 <= or_reduce(nios2_fpu_burst_7_upstream_arb_share_counter_next_value);
  --nios2_fast_fpu/instruction_master nios2_fpu_burst_7/upstream arbiterlock2, which is an e_assign
  nios2_fast_fpu_instruction_master_arbiterlock2 <= nios2_fpu_burst_7_upstream_slavearbiterlockenable2 AND nios2_fast_fpu_instruction_master_continuerequest;
  --nios2_fpu_burst_7_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_fpu_burst_7_upstream_any_continuerequest <= std_logic'('1');
  --nios2_fast_fpu_instruction_master_continuerequest continued request, which is an e_assign
  nios2_fast_fpu_instruction_master_continuerequest <= std_logic'('1');
  internal_nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream <= internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream AND NOT ((nios2_fast_fpu_instruction_master_read AND (((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_instruction_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_instruction_master_latency_counter))))))) OR (nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register)) OR (nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register)))));
  --unique name for nios2_fpu_burst_7_upstream_move_on_to_next_transaction, which is an e_assign
  nios2_fpu_burst_7_upstream_move_on_to_next_transaction <= nios2_fpu_burst_7_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_7_upstream_load_fifo;
  --the currently selected burstcount for nios2_fpu_burst_7_upstream, which is an e_mux
  nios2_fpu_burst_7_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_instruction_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_nios2_fpu_burst_7_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_nios2_fpu_burst_7_upstream : burstcount_fifo_for_nios2_fpu_burst_7_upstream_module
    port map(
      data_out => nios2_fpu_burst_7_upstream_transaction_burst_count,
      empty => nios2_fpu_burst_7_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input42,
      clk => clk,
      data_in => nios2_fpu_burst_7_upstream_selected_burstcount,
      read => nios2_fpu_burst_7_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input43,
      write => module_input44
    );

  module_input42 <= std_logic'('0');
  module_input43 <= std_logic'('0');
  module_input44 <= ((in_a_read_cycle AND NOT nios2_fpu_burst_7_upstream_waits_for_read) AND nios2_fpu_burst_7_upstream_load_fifo) AND NOT ((nios2_fpu_burst_7_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_7_upstream_burstcount_fifo_empty));

  --nios2_fpu_burst_7_upstream current burst minus one, which is an e_assign
  nios2_fpu_burst_7_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_7_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for nios2_fpu_burst_7_upstream, which is an e_mux
  nios2_fpu_burst_7_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_7_upstream_waits_for_read)) AND NOT nios2_fpu_burst_7_upstream_load_fifo))) = '1'), nios2_fpu_burst_7_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_7_upstream_waits_for_read) AND nios2_fpu_burst_7_upstream_this_cycle_is_the_last_burst) AND nios2_fpu_burst_7_upstream_burstcount_fifo_empty))) = '1'), nios2_fpu_burst_7_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((nios2_fpu_burst_7_upstream_this_cycle_is_the_last_burst)) = '1'), nios2_fpu_burst_7_upstream_transaction_burst_count, nios2_fpu_burst_7_upstream_current_burst_minus_one)));
  --the current burst count for nios2_fpu_burst_7_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_7_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((nios2_fpu_burst_7_upstream_readdatavalid_from_sa OR ((NOT nios2_fpu_burst_7_upstream_load_fifo AND ((in_a_read_cycle AND NOT nios2_fpu_burst_7_upstream_waits_for_read)))))) = '1' then 
        nios2_fpu_burst_7_upstream_current_burst <= nios2_fpu_burst_7_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_nios2_fpu_burst_7_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT nios2_fpu_burst_7_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_7_upstream_waits_for_read)) AND nios2_fpu_burst_7_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_7_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_7_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_7_upstream_waits_for_read)) AND NOT nios2_fpu_burst_7_upstream_load_fifo) OR nios2_fpu_burst_7_upstream_this_cycle_is_the_last_burst)) = '1' then 
        nios2_fpu_burst_7_upstream_load_fifo <= p0_nios2_fpu_burst_7_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for nios2_fpu_burst_7_upstream, which is an e_assign
  nios2_fpu_burst_7_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(nios2_fpu_burst_7_upstream_current_burst_minus_one)) AND nios2_fpu_burst_7_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_7_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_7_upstream : rdv_fifo_for_nios2_fast_fpu_instruction_master_to_nios2_fpu_burst_7_upstream_module
    port map(
      data_out => nios2_fast_fpu_instruction_master_rdv_fifo_output_from_nios2_fpu_burst_7_upstream,
      empty => open,
      fifo_contains_ones_n => nios2_fast_fpu_instruction_master_rdv_fifo_empty_nios2_fpu_burst_7_upstream,
      full => open,
      clear_fifo => module_input45,
      clk => clk,
      data_in => internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream,
      read => nios2_fpu_burst_7_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input46,
      write => module_input47
    );

  module_input45 <= std_logic'('0');
  module_input46 <= std_logic'('0');
  module_input47 <= in_a_read_cycle AND NOT nios2_fpu_burst_7_upstream_waits_for_read;

  nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register <= NOT nios2_fast_fpu_instruction_master_rdv_fifo_empty_nios2_fpu_burst_7_upstream;
  --local readdatavalid nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream, which is an e_mux
  nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream <= nios2_fpu_burst_7_upstream_readdatavalid_from_sa;
  --byteaddress mux for nios2_fpu_burst_7/upstream, which is an e_mux
  nios2_fpu_burst_7_upstream_byteaddress <= nios2_fast_fpu_instruction_master_address_to_slave (14 DOWNTO 0);
  --master is always granted when requested
  internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream <= internal_nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream;
  --nios2_fast_fpu/instruction_master saved-grant nios2_fpu_burst_7/upstream, which is an e_assign
  nios2_fast_fpu_instruction_master_saved_grant_nios2_fpu_burst_7_upstream <= internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream;
  --allow new arb cycle for nios2_fpu_burst_7/upstream, which is an e_assign
  nios2_fpu_burst_7_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_fpu_burst_7_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_fpu_burst_7_upstream_master_qreq_vector <= std_logic'('1');
  --nios2_fpu_burst_7_upstream_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_7_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_fpu_burst_7_upstream_begins_xfer) = '1'), nios2_fpu_burst_7_upstream_unreg_firsttransfer, nios2_fpu_burst_7_upstream_reg_firsttransfer);
  --nios2_fpu_burst_7_upstream_unreg_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_7_upstream_unreg_firsttransfer <= NOT ((nios2_fpu_burst_7_upstream_slavearbiterlockenable AND nios2_fpu_burst_7_upstream_any_continuerequest));
  --nios2_fpu_burst_7_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_7_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_7_upstream_begins_xfer) = '1' then 
        nios2_fpu_burst_7_upstream_reg_firsttransfer <= nios2_fpu_burst_7_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_7_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_fpu_burst_7_upstream_beginbursttransfer_internal <= nios2_fpu_burst_7_upstream_begins_xfer;
  --nios2_fpu_burst_7_upstream_read assignment, which is an e_mux
  nios2_fpu_burst_7_upstream_read <= internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream AND nios2_fast_fpu_instruction_master_read;
  --nios2_fpu_burst_7_upstream_write assignment, which is an e_mux
  nios2_fpu_burst_7_upstream_write <= std_logic'('0');
  --nios2_fpu_burst_7_upstream_address mux, which is an e_mux
  nios2_fpu_burst_7_upstream_address <= nios2_fast_fpu_instruction_master_address_to_slave (12 DOWNTO 0);
  --d1_nios2_fpu_burst_7_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_fpu_burst_7_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_fpu_burst_7_upstream_end_xfer <= nios2_fpu_burst_7_upstream_end_xfer;
    end if;

  end process;

  --nios2_fpu_burst_7_upstream_waits_for_read in a cycle, which is an e_mux
  nios2_fpu_burst_7_upstream_waits_for_read <= nios2_fpu_burst_7_upstream_in_a_read_cycle AND internal_nios2_fpu_burst_7_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_7_upstream_in_a_read_cycle assignment, which is an e_assign
  nios2_fpu_burst_7_upstream_in_a_read_cycle <= internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream AND nios2_fast_fpu_instruction_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_fpu_burst_7_upstream_in_a_read_cycle;
  --nios2_fpu_burst_7_upstream_waits_for_write in a cycle, which is an e_mux
  nios2_fpu_burst_7_upstream_waits_for_write <= nios2_fpu_burst_7_upstream_in_a_write_cycle AND internal_nios2_fpu_burst_7_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_7_upstream_in_a_write_cycle assignment, which is an e_assign
  nios2_fpu_burst_7_upstream_in_a_write_cycle <= std_logic'('0');
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_fpu_burst_7_upstream_in_a_write_cycle;
  wait_for_nios2_fpu_burst_7_upstream_counter <= std_logic'('0');
  --nios2_fpu_burst_7_upstream_byteenable byte enable port mux, which is an e_mux
  nios2_fpu_burst_7_upstream_byteenable <= A_EXT (-SIGNED(std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  nios2_fpu_burst_7_upstream_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream <= internal_nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream;
  --vhdl renameroo for output signals
  nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream <= internal_nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream;
  --vhdl renameroo for output signals
  nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream <= internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream;
  --vhdl renameroo for output signals
  nios2_fpu_burst_7_upstream_waitrequest_from_sa <= internal_nios2_fpu_burst_7_upstream_waitrequest_from_sa;
--synthesis translate_off
    --nios2_fpu_burst_7/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --nios2_fast_fpu/instruction_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line75 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_instruction_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line75, now);
          write(write_line75, string'(": "));
          write(write_line75, string'("nios2_fast_fpu/instruction_master drove 0 on its 'burstcount' port while accessing slave nios2_fpu_burst_7/upstream"));
          write(output, write_line75.all);
          deallocate (write_line75);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_7_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_ipl_memory_s1_end_xfer : IN STD_LOGIC;
                 signal ipl_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_7_downstream_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_burst_7_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_7_downstream_granted_ipl_memory_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_requests_ipl_memory_s1 : IN STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_fpu_burst_7_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_burst_7_downstream_latency_counter : OUT STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_7_downstream_readdatavalid : OUT STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_reset_n : OUT STD_LOGIC;
                 signal nios2_fpu_burst_7_downstream_waitrequest : OUT STD_LOGIC
              );
end entity nios2_fpu_burst_7_downstream_arbitrator;


architecture europa of nios2_fpu_burst_7_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_fpu_burst_7_downstream_address_to_slave :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal internal_nios2_fpu_burst_7_downstream_latency_counter :  STD_LOGIC;
                signal internal_nios2_fpu_burst_7_downstream_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_address_last_time :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_7_downstream_burstcount_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_7_downstream_is_granted_some_slave :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_read_but_no_slave_selected :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_read_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_run :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_write_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_nios2_fpu_burst_7_downstream_latency_counter :  STD_LOGIC;
                signal pre_flush_nios2_fpu_burst_7_downstream_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1 OR NOT nios2_fpu_burst_7_downstream_requests_ipl_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_7_downstream_granted_ipl_memory_s1 OR NOT nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1 OR NOT ((nios2_fpu_burst_7_downstream_read OR nios2_fpu_burst_7_downstream_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_7_downstream_read OR nios2_fpu_burst_7_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1 OR NOT ((nios2_fpu_burst_7_downstream_read OR nios2_fpu_burst_7_downstream_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_7_downstream_read OR nios2_fpu_burst_7_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_fpu_burst_7_downstream_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_fpu_burst_7_downstream_address_to_slave <= nios2_fpu_burst_7_downstream_address;
  --nios2_fpu_burst_7_downstream_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_7_downstream_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      nios2_fpu_burst_7_downstream_read_but_no_slave_selected <= (nios2_fpu_burst_7_downstream_read AND nios2_fpu_burst_7_downstream_run) AND NOT nios2_fpu_burst_7_downstream_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  nios2_fpu_burst_7_downstream_is_granted_some_slave <= nios2_fpu_burst_7_downstream_granted_ipl_memory_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_nios2_fpu_burst_7_downstream_readdatavalid <= nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  nios2_fpu_burst_7_downstream_readdatavalid <= nios2_fpu_burst_7_downstream_read_but_no_slave_selected OR pre_flush_nios2_fpu_burst_7_downstream_readdatavalid;
  --nios2_fpu_burst_7/downstream readdata mux, which is an e_mux
  nios2_fpu_burst_7_downstream_readdata <= ipl_memory_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_fpu_burst_7_downstream_waitrequest <= NOT nios2_fpu_burst_7_downstream_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_nios2_fpu_burst_7_downstream_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_nios2_fpu_burst_7_downstream_latency_counter <= p1_nios2_fpu_burst_7_downstream_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_nios2_fpu_burst_7_downstream_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((nios2_fpu_burst_7_downstream_run AND nios2_fpu_burst_7_downstream_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_7_downstream_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_7_downstream_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_7_downstream_requests_ipl_memory_s1))) AND std_logic_vector'("00000000000000000000000000000001")));
  --nios2_fpu_burst_7_downstream_reset_n assignment, which is an e_assign
  nios2_fpu_burst_7_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_fpu_burst_7_downstream_address_to_slave <= internal_nios2_fpu_burst_7_downstream_address_to_slave;
  --vhdl renameroo for output signals
  nios2_fpu_burst_7_downstream_latency_counter <= internal_nios2_fpu_burst_7_downstream_latency_counter;
  --vhdl renameroo for output signals
  nios2_fpu_burst_7_downstream_waitrequest <= internal_nios2_fpu_burst_7_downstream_waitrequest;
--synthesis translate_off
    --nios2_fpu_burst_7_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_7_downstream_address_last_time <= std_logic_vector'("0000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_7_downstream_address_last_time <= nios2_fpu_burst_7_downstream_address;
      end if;

    end process;

    --nios2_fpu_burst_7/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_fpu_burst_7_downstream_waitrequest AND ((nios2_fpu_burst_7_downstream_read OR nios2_fpu_burst_7_downstream_write));
      end if;

    end process;

    --nios2_fpu_burst_7_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line76 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_7_downstream_address /= nios2_fpu_burst_7_downstream_address_last_time))))) = '1' then 
          write(write_line76, now);
          write(write_line76, string'(": "));
          write(write_line76, string'("nios2_fpu_burst_7_downstream_address did not heed wait!!!"));
          write(output, write_line76.all);
          deallocate (write_line76);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_7_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_7_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_7_downstream_burstcount_last_time <= nios2_fpu_burst_7_downstream_burstcount;
      end if;

    end process;

    --nios2_fpu_burst_7_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line77 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_7_downstream_burstcount) /= std_logic'(nios2_fpu_burst_7_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line77, now);
          write(write_line77, string'(": "));
          write(write_line77, string'("nios2_fpu_burst_7_downstream_burstcount did not heed wait!!!"));
          write(output, write_line77.all);
          deallocate (write_line77);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_7_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_7_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_7_downstream_byteenable_last_time <= nios2_fpu_burst_7_downstream_byteenable;
      end if;

    end process;

    --nios2_fpu_burst_7_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line78 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_7_downstream_byteenable /= nios2_fpu_burst_7_downstream_byteenable_last_time))))) = '1' then 
          write(write_line78, now);
          write(write_line78, string'(": "));
          write(write_line78, string'("nios2_fpu_burst_7_downstream_byteenable did not heed wait!!!"));
          write(output, write_line78.all);
          deallocate (write_line78);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_7_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_7_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_7_downstream_read_last_time <= nios2_fpu_burst_7_downstream_read;
      end if;

    end process;

    --nios2_fpu_burst_7_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line79 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_7_downstream_read) /= std_logic'(nios2_fpu_burst_7_downstream_read_last_time)))))) = '1' then 
          write(write_line79, now);
          write(write_line79, string'(": "));
          write(write_line79, string'("nios2_fpu_burst_7_downstream_read did not heed wait!!!"));
          write(output, write_line79.all);
          deallocate (write_line79);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_7_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_7_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_7_downstream_write_last_time <= nios2_fpu_burst_7_downstream_write;
      end if;

    end process;

    --nios2_fpu_burst_7_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line80 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_7_downstream_write) /= std_logic'(nios2_fpu_burst_7_downstream_write_last_time)))))) = '1' then 
          write(write_line80, now);
          write(write_line80, string'(": "));
          write(write_line80, string'("nios2_fpu_burst_7_downstream_write did not heed wait!!!"));
          write(output, write_line80.all);
          deallocate (write_line80);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_7_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_7_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_7_downstream_writedata_last_time <= nios2_fpu_burst_7_downstream_writedata;
      end if;

    end process;

    --nios2_fpu_burst_7_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line81 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_7_downstream_writedata /= nios2_fpu_burst_7_downstream_writedata_last_time)))) AND nios2_fpu_burst_7_downstream_write)) = '1' then 
          write(write_line81, now);
          write(write_line81, string'(": "));
          write(write_line81, string'("nios2_fpu_burst_7_downstream_writedata did not heed wait!!!"));
          write(output, write_line81.all);
          deallocate (write_line81);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity burstcount_fifo_for_nios2_fpu_burst_8_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity burstcount_fifo_for_nios2_fpu_burst_8_upstream_module;


architecture europa of burstcount_fifo_for_nios2_fpu_burst_8_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_2;
  empty <= NOT(full_0);
  full_3 <= std_logic'('0');
  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("0000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("0000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("0000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_8_upstream_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_8_upstream_module;


architecture europa of rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_8_upstream_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_2;
  empty <= NOT(full_0);
  full_3 <= std_logic'('0');
  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_8_upstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fast_fpu_data_master_debugaccess : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_latency_counter : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_write : IN STD_LOGIC;
                 signal nios2_fast_fpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_8_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_8_upstream_readdatavalid : IN STD_LOGIC;
                 signal nios2_fpu_burst_8_upstream_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_nios2_fpu_burst_8_upstream_end_xfer : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register : OUT STD_LOGIC;
                 signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream : OUT STD_LOGIC;
                 signal nios2_fpu_burst_8_upstream_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_burst_8_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_8_upstream_byteaddress : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                 signal nios2_fpu_burst_8_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_8_upstream_debugaccess : OUT STD_LOGIC;
                 signal nios2_fpu_burst_8_upstream_read : OUT STD_LOGIC;
                 signal nios2_fpu_burst_8_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_8_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_fpu_burst_8_upstream_write : OUT STD_LOGIC;
                 signal nios2_fpu_burst_8_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity nios2_fpu_burst_8_upstream_arbitrator;


architecture europa of nios2_fpu_burst_8_upstream_arbitrator is
component burstcount_fifo_for_nios2_fpu_burst_8_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component burstcount_fifo_for_nios2_fpu_burst_8_upstream_module;

component rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_8_upstream_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_8_upstream_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_fpu_burst_8_upstream :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream :  STD_LOGIC;
                signal internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream :  STD_LOGIC;
                signal internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream :  STD_LOGIC;
                signal internal_nios2_fpu_burst_8_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_nios2_fpu_burst_8_upstream_read :  STD_LOGIC;
                signal internal_nios2_fpu_burst_8_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal internal_nios2_fpu_burst_8_upstream_write :  STD_LOGIC;
                signal module_input48 :  STD_LOGIC;
                signal module_input49 :  STD_LOGIC;
                signal module_input50 :  STD_LOGIC;
                signal module_input51 :  STD_LOGIC;
                signal module_input52 :  STD_LOGIC;
                signal module_input53 :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_arbiterlock :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_continuerequest :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_rdv_fifo_empty_nios2_fpu_burst_8_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_rdv_fifo_output_from_nios2_fpu_burst_8_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_saved_grant_nios2_fpu_burst_8_upstream :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_allgrants :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_any_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_arb_counter_enable :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_arb_share_counter :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_arb_share_counter_next_value :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_arb_share_set_values :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_bbt_burstcounter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_begins_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_burstcount_fifo_empty :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_current_burst :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_current_burst_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_end_xfer :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_grant_vector :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_in_a_read_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_in_a_write_cycle :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_load_fifo :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_master_qreq_vector :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_move_on_to_next_transaction :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_next_bbt_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_next_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_readdatavalid_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_reg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_selected_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_this_cycle_is_the_last_burst :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_transaction_burst_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_waits_for_read :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_waits_for_write :  STD_LOGIC;
                signal p0_nios2_fpu_burst_8_upstream_load_fifo :  STD_LOGIC;
                signal wait_for_nios2_fpu_burst_8_upstream_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_fpu_burst_8_upstream_end_xfer;
    end if;

  end process;

  nios2_fpu_burst_8_upstream_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream);
  --assign nios2_fpu_burst_8_upstream_readdatavalid_from_sa = nios2_fpu_burst_8_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_8_upstream_readdatavalid_from_sa <= nios2_fpu_burst_8_upstream_readdatavalid;
  --assign nios2_fpu_burst_8_upstream_readdata_from_sa = nios2_fpu_burst_8_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_burst_8_upstream_readdata_from_sa <= nios2_fpu_burst_8_upstream_readdata;
  internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream <= to_std_logic(((Std_Logic_Vector'(nios2_fast_fpu_data_master_address_to_slave(28 DOWNTO 13) & std_logic_vector'("0000000000000")) = std_logic_vector'("10000000000000000000000000000")))) AND ((nios2_fast_fpu_data_master_read OR nios2_fast_fpu_data_master_write));
  --assign nios2_fpu_burst_8_upstream_waitrequest_from_sa = nios2_fpu_burst_8_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_fpu_burst_8_upstream_waitrequest_from_sa <= nios2_fpu_burst_8_upstream_waitrequest;
  --nios2_fpu_burst_8_upstream_arb_share_counter set values, which is an e_mux
  nios2_fpu_burst_8_upstream_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream)) = '1'), (A_WE_StdLogicVector((std_logic'((nios2_fast_fpu_data_master_write)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001"))), std_logic_vector'("00000000000000000000000000000001")), 6);
  --nios2_fpu_burst_8_upstream_non_bursting_master_requests mux, which is an e_mux
  nios2_fpu_burst_8_upstream_non_bursting_master_requests <= std_logic'('0');
  --nios2_fpu_burst_8_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_fpu_burst_8_upstream_any_bursting_master_saved_grant <= nios2_fast_fpu_data_master_saved_grant_nios2_fpu_burst_8_upstream;
  --nios2_fpu_burst_8_upstream_arb_share_counter_next_value assignment, which is an e_assign
  nios2_fpu_burst_8_upstream_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_8_upstream_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_8_upstream_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_fpu_burst_8_upstream_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_8_upstream_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 6);
  --nios2_fpu_burst_8_upstream_allgrants all slave grants, which is an e_mux
  nios2_fpu_burst_8_upstream_allgrants <= nios2_fpu_burst_8_upstream_grant_vector;
  --nios2_fpu_burst_8_upstream_end_xfer assignment, which is an e_assign
  nios2_fpu_burst_8_upstream_end_xfer <= NOT ((nios2_fpu_burst_8_upstream_waits_for_read OR nios2_fpu_burst_8_upstream_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_fpu_burst_8_upstream arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_fpu_burst_8_upstream <= nios2_fpu_burst_8_upstream_end_xfer AND (((NOT nios2_fpu_burst_8_upstream_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_fpu_burst_8_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_fpu_burst_8_upstream_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_fpu_burst_8_upstream AND nios2_fpu_burst_8_upstream_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_8_upstream AND NOT nios2_fpu_burst_8_upstream_non_bursting_master_requests));
  --nios2_fpu_burst_8_upstream_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_8_upstream_arb_share_counter <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_8_upstream_arb_counter_enable) = '1' then 
        nios2_fpu_burst_8_upstream_arb_share_counter <= nios2_fpu_burst_8_upstream_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_8_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_8_upstream_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_fpu_burst_8_upstream_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_fpu_burst_8_upstream)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_burst_8_upstream AND NOT nios2_fpu_burst_8_upstream_non_bursting_master_requests)))) = '1' then 
        nios2_fpu_burst_8_upstream_slavearbiterlockenable <= or_reduce(nios2_fpu_burst_8_upstream_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --nios2_fast_fpu/data_master nios2_fpu_burst_8/upstream arbiterlock, which is an e_assign
  nios2_fast_fpu_data_master_arbiterlock <= nios2_fpu_burst_8_upstream_slavearbiterlockenable AND nios2_fast_fpu_data_master_continuerequest;
  --nios2_fpu_burst_8_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_fpu_burst_8_upstream_slavearbiterlockenable2 <= or_reduce(nios2_fpu_burst_8_upstream_arb_share_counter_next_value);
  --nios2_fast_fpu/data_master nios2_fpu_burst_8/upstream arbiterlock2, which is an e_assign
  nios2_fast_fpu_data_master_arbiterlock2 <= nios2_fpu_burst_8_upstream_slavearbiterlockenable2 AND nios2_fast_fpu_data_master_continuerequest;
  --nios2_fpu_burst_8_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_fpu_burst_8_upstream_any_continuerequest <= std_logic'('1');
  --nios2_fast_fpu_data_master_continuerequest continued request, which is an e_assign
  nios2_fast_fpu_data_master_continuerequest <= std_logic'('1');
  internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream <= internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream AND NOT ((nios2_fast_fpu_data_master_read AND ((((to_std_logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_data_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_data_master_latency_counter))))))) OR (nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register)) OR (nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register)) OR (nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register)))));
  --unique name for nios2_fpu_burst_8_upstream_move_on_to_next_transaction, which is an e_assign
  nios2_fpu_burst_8_upstream_move_on_to_next_transaction <= nios2_fpu_burst_8_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_8_upstream_load_fifo;
  --the currently selected burstcount for nios2_fpu_burst_8_upstream, which is an e_mux
  nios2_fpu_burst_8_upstream_selected_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --burstcount_fifo_for_nios2_fpu_burst_8_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_nios2_fpu_burst_8_upstream : burstcount_fifo_for_nios2_fpu_burst_8_upstream_module
    port map(
      data_out => nios2_fpu_burst_8_upstream_transaction_burst_count,
      empty => nios2_fpu_burst_8_upstream_burstcount_fifo_empty,
      fifo_contains_ones_n => open,
      full => open,
      clear_fifo => module_input48,
      clk => clk,
      data_in => nios2_fpu_burst_8_upstream_selected_burstcount,
      read => nios2_fpu_burst_8_upstream_this_cycle_is_the_last_burst,
      reset_n => reset_n,
      sync_reset => module_input49,
      write => module_input50
    );

  module_input48 <= std_logic'('0');
  module_input49 <= std_logic'('0');
  module_input50 <= ((in_a_read_cycle AND NOT nios2_fpu_burst_8_upstream_waits_for_read) AND nios2_fpu_burst_8_upstream_load_fifo) AND NOT ((nios2_fpu_burst_8_upstream_this_cycle_is_the_last_burst AND nios2_fpu_burst_8_upstream_burstcount_fifo_empty));

  --nios2_fpu_burst_8_upstream current burst minus one, which is an e_assign
  nios2_fpu_burst_8_upstream_current_burst_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_8_upstream_current_burst)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --what to load in current_burst, for nios2_fpu_burst_8_upstream, which is an e_mux
  nios2_fpu_burst_8_upstream_next_burst_count <= A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_8_upstream_waits_for_read)) AND NOT nios2_fpu_burst_8_upstream_load_fifo))) = '1'), nios2_fpu_burst_8_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_8_upstream_waits_for_read) AND nios2_fpu_burst_8_upstream_this_cycle_is_the_last_burst) AND nios2_fpu_burst_8_upstream_burstcount_fifo_empty))) = '1'), nios2_fpu_burst_8_upstream_selected_burstcount, A_WE_StdLogicVector((std_logic'((nios2_fpu_burst_8_upstream_this_cycle_is_the_last_burst)) = '1'), nios2_fpu_burst_8_upstream_transaction_burst_count, nios2_fpu_burst_8_upstream_current_burst_minus_one)));
  --the current burst count for nios2_fpu_burst_8_upstream, to be decremented, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_8_upstream_current_burst <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((nios2_fpu_burst_8_upstream_readdatavalid_from_sa OR ((NOT nios2_fpu_burst_8_upstream_load_fifo AND ((in_a_read_cycle AND NOT nios2_fpu_burst_8_upstream_waits_for_read)))))) = '1' then 
        nios2_fpu_burst_8_upstream_current_burst <= nios2_fpu_burst_8_upstream_next_burst_count;
      end if;
    end if;

  end process;

  --a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  p0_nios2_fpu_burst_8_upstream_load_fifo <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((NOT nios2_fpu_burst_8_upstream_load_fifo)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_8_upstream_waits_for_read)) AND nios2_fpu_burst_8_upstream_load_fifo))) = '1'), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_8_upstream_burstcount_fifo_empty))))));
  --whether to load directly to the counter or to the fifo, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_8_upstream_load_fifo <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((((in_a_read_cycle AND NOT nios2_fpu_burst_8_upstream_waits_for_read)) AND NOT nios2_fpu_burst_8_upstream_load_fifo) OR nios2_fpu_burst_8_upstream_this_cycle_is_the_last_burst)) = '1' then 
        nios2_fpu_burst_8_upstream_load_fifo <= p0_nios2_fpu_burst_8_upstream_load_fifo;
      end if;
    end if;

  end process;

  --the last cycle in the burst for nios2_fpu_burst_8_upstream, which is an e_assign
  nios2_fpu_burst_8_upstream_this_cycle_is_the_last_burst <= NOT (or_reduce(nios2_fpu_burst_8_upstream_current_burst_minus_one)) AND nios2_fpu_burst_8_upstream_readdatavalid_from_sa;
  --rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_8_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_8_upstream : rdv_fifo_for_nios2_fast_fpu_data_master_to_nios2_fpu_burst_8_upstream_module
    port map(
      data_out => nios2_fast_fpu_data_master_rdv_fifo_output_from_nios2_fpu_burst_8_upstream,
      empty => open,
      fifo_contains_ones_n => nios2_fast_fpu_data_master_rdv_fifo_empty_nios2_fpu_burst_8_upstream,
      full => open,
      clear_fifo => module_input51,
      clk => clk,
      data_in => internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream,
      read => nios2_fpu_burst_8_upstream_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input52,
      write => module_input53
    );

  module_input51 <= std_logic'('0');
  module_input52 <= std_logic'('0');
  module_input53 <= in_a_read_cycle AND NOT nios2_fpu_burst_8_upstream_waits_for_read;

  nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register <= NOT nios2_fast_fpu_data_master_rdv_fifo_empty_nios2_fpu_burst_8_upstream;
  --local readdatavalid nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream, which is an e_mux
  nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream <= nios2_fpu_burst_8_upstream_readdatavalid_from_sa;
  --nios2_fpu_burst_8_upstream_writedata mux, which is an e_mux
  nios2_fpu_burst_8_upstream_writedata <= nios2_fast_fpu_data_master_writedata;
  --byteaddress mux for nios2_fpu_burst_8/upstream, which is an e_mux
  nios2_fpu_burst_8_upstream_byteaddress <= nios2_fast_fpu_data_master_address_to_slave (14 DOWNTO 0);
  --master is always granted when requested
  internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream <= internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream;
  --nios2_fast_fpu/data_master saved-grant nios2_fpu_burst_8/upstream, which is an e_assign
  nios2_fast_fpu_data_master_saved_grant_nios2_fpu_burst_8_upstream <= internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream;
  --allow new arb cycle for nios2_fpu_burst_8/upstream, which is an e_assign
  nios2_fpu_burst_8_upstream_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_fpu_burst_8_upstream_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_fpu_burst_8_upstream_master_qreq_vector <= std_logic'('1');
  --nios2_fpu_burst_8_upstream_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_8_upstream_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_fpu_burst_8_upstream_begins_xfer) = '1'), nios2_fpu_burst_8_upstream_unreg_firsttransfer, nios2_fpu_burst_8_upstream_reg_firsttransfer);
  --nios2_fpu_burst_8_upstream_unreg_firsttransfer first transaction, which is an e_assign
  nios2_fpu_burst_8_upstream_unreg_firsttransfer <= NOT ((nios2_fpu_burst_8_upstream_slavearbiterlockenable AND nios2_fpu_burst_8_upstream_any_continuerequest));
  --nios2_fpu_burst_8_upstream_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_8_upstream_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_8_upstream_begins_xfer) = '1' then 
        nios2_fpu_burst_8_upstream_reg_firsttransfer <= nios2_fpu_burst_8_upstream_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_8_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  nios2_fpu_burst_8_upstream_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_nios2_fpu_burst_8_upstream_write) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_8_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (internal_nios2_fpu_burst_8_upstream_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_nios2_fpu_burst_8_upstream_read) AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_8_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("000000000000000000000000000000") & (nios2_fpu_burst_8_upstream_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 3);
  --nios2_fpu_burst_8_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_burst_8_upstream_bbt_burstcounter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_burst_8_upstream_begins_xfer) = '1' then 
        nios2_fpu_burst_8_upstream_bbt_burstcounter <= nios2_fpu_burst_8_upstream_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --nios2_fpu_burst_8_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_fpu_burst_8_upstream_beginbursttransfer_internal <= nios2_fpu_burst_8_upstream_begins_xfer AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_8_upstream_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --nios2_fpu_burst_8_upstream_read assignment, which is an e_mux
  internal_nios2_fpu_burst_8_upstream_read <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream AND nios2_fast_fpu_data_master_read;
  --nios2_fpu_burst_8_upstream_write assignment, which is an e_mux
  internal_nios2_fpu_burst_8_upstream_write <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream AND nios2_fast_fpu_data_master_write;
  --nios2_fpu_burst_8_upstream_address mux, which is an e_mux
  nios2_fpu_burst_8_upstream_address <= nios2_fast_fpu_data_master_address_to_slave (12 DOWNTO 0);
  --d1_nios2_fpu_burst_8_upstream_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_fpu_burst_8_upstream_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_fpu_burst_8_upstream_end_xfer <= nios2_fpu_burst_8_upstream_end_xfer;
    end if;

  end process;

  --nios2_fpu_burst_8_upstream_waits_for_read in a cycle, which is an e_mux
  nios2_fpu_burst_8_upstream_waits_for_read <= nios2_fpu_burst_8_upstream_in_a_read_cycle AND internal_nios2_fpu_burst_8_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_8_upstream_in_a_read_cycle assignment, which is an e_assign
  nios2_fpu_burst_8_upstream_in_a_read_cycle <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream AND nios2_fast_fpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_fpu_burst_8_upstream_in_a_read_cycle;
  --nios2_fpu_burst_8_upstream_waits_for_write in a cycle, which is an e_mux
  nios2_fpu_burst_8_upstream_waits_for_write <= nios2_fpu_burst_8_upstream_in_a_write_cycle AND internal_nios2_fpu_burst_8_upstream_waitrequest_from_sa;
  --nios2_fpu_burst_8_upstream_in_a_write_cycle assignment, which is an e_assign
  nios2_fpu_burst_8_upstream_in_a_write_cycle <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream AND nios2_fast_fpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_fpu_burst_8_upstream_in_a_write_cycle;
  wait_for_nios2_fpu_burst_8_upstream_counter <= std_logic'('0');
  --nios2_fpu_burst_8_upstream_byteenable byte enable port mux, which is an e_mux
  nios2_fpu_burst_8_upstream_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --burstcount mux, which is an e_mux
  internal_nios2_fpu_burst_8_upstream_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_burstcount)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --debugaccess mux, which is an e_mux
  nios2_fpu_burst_8_upstream_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream <= internal_nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream;
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream <= internal_nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream;
  --vhdl renameroo for output signals
  nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream <= internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream;
  --vhdl renameroo for output signals
  nios2_fpu_burst_8_upstream_burstcount <= internal_nios2_fpu_burst_8_upstream_burstcount;
  --vhdl renameroo for output signals
  nios2_fpu_burst_8_upstream_read <= internal_nios2_fpu_burst_8_upstream_read;
  --vhdl renameroo for output signals
  nios2_fpu_burst_8_upstream_waitrequest_from_sa <= internal_nios2_fpu_burst_8_upstream_waitrequest_from_sa;
  --vhdl renameroo for output signals
  nios2_fpu_burst_8_upstream_write <= internal_nios2_fpu_burst_8_upstream_write;
--synthesis translate_off
    --nios2_fpu_burst_8/upstream enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --nios2_fast_fpu/data_master non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line82 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (nios2_fast_fpu_data_master_burstcount)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line82, now);
          write(write_line82, string'(": "));
          write(write_line82, string'("nios2_fast_fpu/data_master drove 0 on its 'burstcount' port while accessing slave nios2_fpu_burst_8/upstream"));
          write(output, write_line82.all);
          deallocate (write_line82);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_burst_8_downstream_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_nios2_fpu_clock_0_in_end_xfer : IN STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_burst_8_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in : IN STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in : IN STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_read_data_valid_nios2_fpu_clock_0_in : IN STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in : IN STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_clock_0_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_clock_0_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_fpu_burst_8_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_burst_8_downstream_latency_counter : OUT STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_burst_8_downstream_readdatavalid : OUT STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_reset_n : OUT STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_waitrequest : OUT STD_LOGIC
              );
end entity nios2_fpu_burst_8_downstream_arbitrator;


architecture europa of nios2_fpu_burst_8_downstream_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_fpu_burst_8_downstream_address_to_slave :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal internal_nios2_fpu_burst_8_downstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_address_last_time :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_8_downstream_burstcount_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_8_downstream_read_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_run :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_write_last_time :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pre_flush_nios2_fpu_burst_8_downstream_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in OR NOT nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in OR NOT ((nios2_fpu_burst_8_downstream_read OR nios2_fpu_burst_8_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_clock_0_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_8_downstream_read OR nios2_fpu_burst_8_downstream_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in OR NOT ((nios2_fpu_burst_8_downstream_read OR nios2_fpu_burst_8_downstream_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_clock_0_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_8_downstream_read OR nios2_fpu_burst_8_downstream_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_fpu_burst_8_downstream_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_fpu_burst_8_downstream_address_to_slave <= nios2_fpu_burst_8_downstream_address;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_nios2_fpu_burst_8_downstream_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  nios2_fpu_burst_8_downstream_readdatavalid <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_nios2_fpu_burst_8_downstream_readdatavalid)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_8_downstream_read_data_valid_nios2_fpu_clock_0_in)))));
  --nios2_fpu_burst_8/downstream readdata mux, which is an e_mux
  nios2_fpu_burst_8_downstream_readdata <= nios2_fpu_clock_0_in_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_fpu_burst_8_downstream_waitrequest <= NOT nios2_fpu_burst_8_downstream_run;
  --latent max counter, which is an e_assign
  nios2_fpu_burst_8_downstream_latency_counter <= std_logic'('0');
  --nios2_fpu_burst_8_downstream_reset_n assignment, which is an e_assign
  nios2_fpu_burst_8_downstream_reset_n <= reset_n;
  --vhdl renameroo for output signals
  nios2_fpu_burst_8_downstream_address_to_slave <= internal_nios2_fpu_burst_8_downstream_address_to_slave;
  --vhdl renameroo for output signals
  nios2_fpu_burst_8_downstream_waitrequest <= internal_nios2_fpu_burst_8_downstream_waitrequest;
--synthesis translate_off
    --nios2_fpu_burst_8_downstream_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_8_downstream_address_last_time <= std_logic_vector'("0000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_8_downstream_address_last_time <= nios2_fpu_burst_8_downstream_address;
      end if;

    end process;

    --nios2_fpu_burst_8/downstream waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_fpu_burst_8_downstream_waitrequest AND ((nios2_fpu_burst_8_downstream_read OR nios2_fpu_burst_8_downstream_write));
      end if;

    end process;

    --nios2_fpu_burst_8_downstream_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line83 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_8_downstream_address /= nios2_fpu_burst_8_downstream_address_last_time))))) = '1' then 
          write(write_line83, now);
          write(write_line83, string'(": "));
          write(write_line83, string'("nios2_fpu_burst_8_downstream_address did not heed wait!!!"));
          write(output, write_line83.all);
          deallocate (write_line83);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_8_downstream_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_8_downstream_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_8_downstream_burstcount_last_time <= nios2_fpu_burst_8_downstream_burstcount;
      end if;

    end process;

    --nios2_fpu_burst_8_downstream_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line84 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_8_downstream_burstcount) /= std_logic'(nios2_fpu_burst_8_downstream_burstcount_last_time)))))) = '1' then 
          write(write_line84, now);
          write(write_line84, string'(": "));
          write(write_line84, string'("nios2_fpu_burst_8_downstream_burstcount did not heed wait!!!"));
          write(output, write_line84.all);
          deallocate (write_line84);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_8_downstream_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_8_downstream_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_8_downstream_byteenable_last_time <= nios2_fpu_burst_8_downstream_byteenable;
      end if;

    end process;

    --nios2_fpu_burst_8_downstream_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line85 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_8_downstream_byteenable /= nios2_fpu_burst_8_downstream_byteenable_last_time))))) = '1' then 
          write(write_line85, now);
          write(write_line85, string'(": "));
          write(write_line85, string'("nios2_fpu_burst_8_downstream_byteenable did not heed wait!!!"));
          write(output, write_line85.all);
          deallocate (write_line85);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_8_downstream_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_8_downstream_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_8_downstream_read_last_time <= nios2_fpu_burst_8_downstream_read;
      end if;

    end process;

    --nios2_fpu_burst_8_downstream_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line86 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_8_downstream_read) /= std_logic'(nios2_fpu_burst_8_downstream_read_last_time)))))) = '1' then 
          write(write_line86, now);
          write(write_line86, string'(": "));
          write(write_line86, string'("nios2_fpu_burst_8_downstream_read did not heed wait!!!"));
          write(output, write_line86.all);
          deallocate (write_line86);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_8_downstream_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_8_downstream_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_8_downstream_write_last_time <= nios2_fpu_burst_8_downstream_write;
      end if;

    end process;

    --nios2_fpu_burst_8_downstream_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line87 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_burst_8_downstream_write) /= std_logic'(nios2_fpu_burst_8_downstream_write_last_time)))))) = '1' then 
          write(write_line87, now);
          write(write_line87, string'(": "));
          write(write_line87, string'("nios2_fpu_burst_8_downstream_write did not heed wait!!!"));
          write(output, write_line87.all);
          deallocate (write_line87);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_8_downstream_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_burst_8_downstream_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_burst_8_downstream_writedata_last_time <= nios2_fpu_burst_8_downstream_writedata;
      end if;

    end process;

    --nios2_fpu_burst_8_downstream_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line88 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_burst_8_downstream_writedata /= nios2_fpu_burst_8_downstream_writedata_last_time)))) AND nios2_fpu_burst_8_downstream_write)) = '1' then 
          write(write_line88, now);
          write(write_line88, string'(": "));
          write(write_line88, string'("nios2_fpu_burst_8_downstream_writedata did not heed wait!!!"));
          write(output, write_line88.all);
          deallocate (write_line88);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_clock_0_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_burst_8_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_8_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_burst_8_downstream_latency_counter : IN STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_nativeaddress : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_burst_8_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_clock_0_in_endofpacket : IN STD_LOGIC;
                 signal nios2_fpu_clock_0_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_clock_0_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_nios2_fpu_clock_0_in_end_xfer : OUT STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in : OUT STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in : OUT STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_read_data_valid_nios2_fpu_clock_0_in : OUT STD_LOGIC;
                 signal nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in : OUT STD_LOGIC;
                 signal nios2_fpu_clock_0_in_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_clock_0_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_clock_0_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal nios2_fpu_clock_0_in_nativeaddress : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal nios2_fpu_clock_0_in_read : OUT STD_LOGIC;
                 signal nios2_fpu_clock_0_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_clock_0_in_reset_n : OUT STD_LOGIC;
                 signal nios2_fpu_clock_0_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal nios2_fpu_clock_0_in_write : OUT STD_LOGIC;
                 signal nios2_fpu_clock_0_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity nios2_fpu_clock_0_in_arbitrator;


architecture europa of nios2_fpu_clock_0_in_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_nios2_fpu_clock_0_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in :  STD_LOGIC;
                signal internal_nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in :  STD_LOGIC;
                signal internal_nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in :  STD_LOGIC;
                signal internal_nios2_fpu_clock_0_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_arbiterlock :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_arbiterlock2 :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_saved_grant_nios2_fpu_clock_0_in :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_allgrants :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_allow_new_arb_cycle :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_any_continuerequest :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_arb_counter_enable :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_arb_share_counter :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_clock_0_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_clock_0_in_arb_share_set_values :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_clock_0_in_beginbursttransfer_internal :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_begins_xfer :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_end_xfer :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_grant_vector :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_in_a_read_cycle :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_in_a_write_cycle :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_master_qreq_vector :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_non_bursting_master_requests :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_reg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_slavearbiterlockenable :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_unreg_firsttransfer :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_waits_for_read :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_waits_for_write :  STD_LOGIC;
                signal wait_for_nios2_fpu_clock_0_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT nios2_fpu_clock_0_in_end_xfer;
    end if;

  end process;

  nios2_fpu_clock_0_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in);
  --assign nios2_fpu_clock_0_in_readdata_from_sa = nios2_fpu_clock_0_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_clock_0_in_readdata_from_sa <= nios2_fpu_clock_0_in_readdata;
  internal_nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_8_downstream_read OR nios2_fpu_burst_8_downstream_write)))))));
  --assign nios2_fpu_clock_0_in_waitrequest_from_sa = nios2_fpu_clock_0_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_nios2_fpu_clock_0_in_waitrequest_from_sa <= nios2_fpu_clock_0_in_waitrequest;
  --nios2_fpu_clock_0_in_arb_share_counter set values, which is an e_mux
  nios2_fpu_clock_0_in_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_8_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001")), 4);
  --nios2_fpu_clock_0_in_non_bursting_master_requests mux, which is an e_mux
  nios2_fpu_clock_0_in_non_bursting_master_requests <= std_logic'('0');
  --nios2_fpu_clock_0_in_any_bursting_master_saved_grant mux, which is an e_mux
  nios2_fpu_clock_0_in_any_bursting_master_saved_grant <= nios2_fpu_burst_8_downstream_saved_grant_nios2_fpu_clock_0_in;
  --nios2_fpu_clock_0_in_arb_share_counter_next_value assignment, which is an e_assign
  nios2_fpu_clock_0_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(nios2_fpu_clock_0_in_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_clock_0_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(nios2_fpu_clock_0_in_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_clock_0_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 4);
  --nios2_fpu_clock_0_in_allgrants all slave grants, which is an e_mux
  nios2_fpu_clock_0_in_allgrants <= nios2_fpu_clock_0_in_grant_vector;
  --nios2_fpu_clock_0_in_end_xfer assignment, which is an e_assign
  nios2_fpu_clock_0_in_end_xfer <= NOT ((nios2_fpu_clock_0_in_waits_for_read OR nios2_fpu_clock_0_in_waits_for_write));
  --end_xfer_arb_share_counter_term_nios2_fpu_clock_0_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_nios2_fpu_clock_0_in <= nios2_fpu_clock_0_in_end_xfer AND (((NOT nios2_fpu_clock_0_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --nios2_fpu_clock_0_in_arb_share_counter arbitration counter enable, which is an e_assign
  nios2_fpu_clock_0_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_nios2_fpu_clock_0_in AND nios2_fpu_clock_0_in_allgrants)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_clock_0_in AND NOT nios2_fpu_clock_0_in_non_bursting_master_requests));
  --nios2_fpu_clock_0_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_clock_0_in_arb_share_counter <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_clock_0_in_arb_counter_enable) = '1' then 
        nios2_fpu_clock_0_in_arb_share_counter <= nios2_fpu_clock_0_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_fpu_clock_0_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_clock_0_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((nios2_fpu_clock_0_in_master_qreq_vector AND end_xfer_arb_share_counter_term_nios2_fpu_clock_0_in)) OR ((end_xfer_arb_share_counter_term_nios2_fpu_clock_0_in AND NOT nios2_fpu_clock_0_in_non_bursting_master_requests)))) = '1' then 
        nios2_fpu_clock_0_in_slavearbiterlockenable <= or_reduce(nios2_fpu_clock_0_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --nios2_fpu_burst_8/downstream nios2_fpu_clock_0/in arbiterlock, which is an e_assign
  nios2_fpu_burst_8_downstream_arbiterlock <= nios2_fpu_clock_0_in_slavearbiterlockenable AND nios2_fpu_burst_8_downstream_continuerequest;
  --nios2_fpu_clock_0_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  nios2_fpu_clock_0_in_slavearbiterlockenable2 <= or_reduce(nios2_fpu_clock_0_in_arb_share_counter_next_value);
  --nios2_fpu_burst_8/downstream nios2_fpu_clock_0/in arbiterlock2, which is an e_assign
  nios2_fpu_burst_8_downstream_arbiterlock2 <= nios2_fpu_clock_0_in_slavearbiterlockenable2 AND nios2_fpu_burst_8_downstream_continuerequest;
  --nios2_fpu_clock_0_in_any_continuerequest at least one master continues requesting, which is an e_assign
  nios2_fpu_clock_0_in_any_continuerequest <= std_logic'('1');
  --nios2_fpu_burst_8_downstream_continuerequest continued request, which is an e_assign
  nios2_fpu_burst_8_downstream_continuerequest <= std_logic'('1');
  internal_nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in <= internal_nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in AND NOT ((nios2_fpu_burst_8_downstream_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_8_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid nios2_fpu_burst_8_downstream_read_data_valid_nios2_fpu_clock_0_in, which is an e_mux
  nios2_fpu_burst_8_downstream_read_data_valid_nios2_fpu_clock_0_in <= (internal_nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in AND nios2_fpu_burst_8_downstream_read) AND NOT nios2_fpu_clock_0_in_waits_for_read;
  --nios2_fpu_clock_0_in_writedata mux, which is an e_mux
  nios2_fpu_clock_0_in_writedata <= nios2_fpu_burst_8_downstream_writedata;
  --assign nios2_fpu_clock_0_in_endofpacket_from_sa = nios2_fpu_clock_0_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  nios2_fpu_clock_0_in_endofpacket_from_sa <= nios2_fpu_clock_0_in_endofpacket;
  --master is always granted when requested
  internal_nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in <= internal_nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in;
  --nios2_fpu_burst_8/downstream saved-grant nios2_fpu_clock_0/in, which is an e_assign
  nios2_fpu_burst_8_downstream_saved_grant_nios2_fpu_clock_0_in <= internal_nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in;
  --allow new arb cycle for nios2_fpu_clock_0/in, which is an e_assign
  nios2_fpu_clock_0_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  nios2_fpu_clock_0_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  nios2_fpu_clock_0_in_master_qreq_vector <= std_logic'('1');
  --nios2_fpu_clock_0_in_reset_n assignment, which is an e_assign
  nios2_fpu_clock_0_in_reset_n <= reset_n;
  --nios2_fpu_clock_0_in_firsttransfer first transaction, which is an e_assign
  nios2_fpu_clock_0_in_firsttransfer <= A_WE_StdLogic((std_logic'(nios2_fpu_clock_0_in_begins_xfer) = '1'), nios2_fpu_clock_0_in_unreg_firsttransfer, nios2_fpu_clock_0_in_reg_firsttransfer);
  --nios2_fpu_clock_0_in_unreg_firsttransfer first transaction, which is an e_assign
  nios2_fpu_clock_0_in_unreg_firsttransfer <= NOT ((nios2_fpu_clock_0_in_slavearbiterlockenable AND nios2_fpu_clock_0_in_any_continuerequest));
  --nios2_fpu_clock_0_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      nios2_fpu_clock_0_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(nios2_fpu_clock_0_in_begins_xfer) = '1' then 
        nios2_fpu_clock_0_in_reg_firsttransfer <= nios2_fpu_clock_0_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --nios2_fpu_clock_0_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  nios2_fpu_clock_0_in_beginbursttransfer_internal <= nios2_fpu_clock_0_in_begins_xfer;
  --nios2_fpu_clock_0_in_read assignment, which is an e_mux
  nios2_fpu_clock_0_in_read <= internal_nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in AND nios2_fpu_burst_8_downstream_read;
  --nios2_fpu_clock_0_in_write assignment, which is an e_mux
  nios2_fpu_clock_0_in_write <= internal_nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in AND nios2_fpu_burst_8_downstream_write;
  --nios2_fpu_clock_0_in_address mux, which is an e_mux
  nios2_fpu_clock_0_in_address <= nios2_fpu_burst_8_downstream_address_to_slave;
  --slaveid nios2_fpu_clock_0_in_nativeaddress nativeaddress mux, which is an e_mux
  nios2_fpu_clock_0_in_nativeaddress <= nios2_fpu_burst_8_downstream_nativeaddress (10 DOWNTO 0);
  --d1_nios2_fpu_clock_0_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_nios2_fpu_clock_0_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_nios2_fpu_clock_0_in_end_xfer <= nios2_fpu_clock_0_in_end_xfer;
    end if;

  end process;

  --nios2_fpu_clock_0_in_waits_for_read in a cycle, which is an e_mux
  nios2_fpu_clock_0_in_waits_for_read <= nios2_fpu_clock_0_in_in_a_read_cycle AND internal_nios2_fpu_clock_0_in_waitrequest_from_sa;
  --nios2_fpu_clock_0_in_in_a_read_cycle assignment, which is an e_assign
  nios2_fpu_clock_0_in_in_a_read_cycle <= internal_nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in AND nios2_fpu_burst_8_downstream_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= nios2_fpu_clock_0_in_in_a_read_cycle;
  --nios2_fpu_clock_0_in_waits_for_write in a cycle, which is an e_mux
  nios2_fpu_clock_0_in_waits_for_write <= nios2_fpu_clock_0_in_in_a_write_cycle AND internal_nios2_fpu_clock_0_in_waitrequest_from_sa;
  --nios2_fpu_clock_0_in_in_a_write_cycle assignment, which is an e_assign
  nios2_fpu_clock_0_in_in_a_write_cycle <= internal_nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in AND nios2_fpu_burst_8_downstream_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= nios2_fpu_clock_0_in_in_a_write_cycle;
  wait_for_nios2_fpu_clock_0_in_counter <= std_logic'('0');
  --nios2_fpu_clock_0_in_byteenable byte enable port mux, which is an e_mux
  nios2_fpu_clock_0_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_8_downstream_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in <= internal_nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in;
  --vhdl renameroo for output signals
  nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in <= internal_nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in;
  --vhdl renameroo for output signals
  nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in <= internal_nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in;
  --vhdl renameroo for output signals
  nios2_fpu_clock_0_in_waitrequest_from_sa <= internal_nios2_fpu_clock_0_in_waitrequest_from_sa;
--synthesis translate_off
    --nios2_fpu_clock_0/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --nios2_fpu_burst_8/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line89 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_burst_8_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line89, now);
          write(write_line89, string'(": "));
          write(write_line89, string'("nios2_fpu_burst_8/downstream drove 0 on its 'arbitrationshare' port while accessing slave nios2_fpu_clock_0/in"));
          write(output, write_line89.all);
          deallocate (write_line89);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_8/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line90 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_8_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line90, now);
          write(write_line90, string'(": "));
          write(write_line90, string'("nios2_fpu_burst_8/downstream drove 0 on its 'burstcount' port while accessing slave nios2_fpu_clock_0/in"));
          write(output, write_line90.all);
          deallocate (write_line90);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity nios2_fpu_clock_0_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_peripheral_bridge_s1_end_xfer : IN STD_LOGIC;
                 signal nios2_fpu_clock_0_out_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_clock_0_out_granted_peripheral_bridge_s1 : IN STD_LOGIC;
                 signal nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1 : IN STD_LOGIC;
                 signal nios2_fpu_clock_0_out_read : IN STD_LOGIC;
                 signal nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1 : IN STD_LOGIC;
                 signal nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1_shift_register : IN STD_LOGIC;
                 signal nios2_fpu_clock_0_out_requests_peripheral_bridge_s1 : IN STD_LOGIC;
                 signal nios2_fpu_clock_0_out_write : IN STD_LOGIC;
                 signal nios2_fpu_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal peripheral_bridge_s1_endofpacket_from_sa : IN STD_LOGIC;
                 signal peripheral_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal peripheral_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal nios2_fpu_clock_0_out_address_to_slave : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_clock_0_out_endofpacket : OUT STD_LOGIC;
                 signal nios2_fpu_clock_0_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal nios2_fpu_clock_0_out_reset_n : OUT STD_LOGIC;
                 signal nios2_fpu_clock_0_out_waitrequest : OUT STD_LOGIC
              );
end entity nios2_fpu_clock_0_out_arbitrator;


architecture europa of nios2_fpu_clock_0_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_nios2_fpu_clock_0_out_address_to_slave :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal internal_nios2_fpu_clock_0_out_waitrequest :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_address_last_time :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_clock_0_out_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_clock_0_out_read_last_time :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_run :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_write_last_time :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_1 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1 OR nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1) OR NOT nios2_fpu_clock_0_out_requests_peripheral_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1 OR NOT nios2_fpu_clock_0_out_read) OR ((nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1 AND nios2_fpu_clock_0_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1 OR NOT ((nios2_fpu_clock_0_out_read OR nios2_fpu_clock_0_out_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT peripheral_bridge_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_clock_0_out_read OR nios2_fpu_clock_0_out_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  nios2_fpu_clock_0_out_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_nios2_fpu_clock_0_out_address_to_slave <= nios2_fpu_clock_0_out_address;
  --nios2_fpu_clock_0/out readdata mux, which is an e_mux
  nios2_fpu_clock_0_out_readdata <= peripheral_bridge_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_nios2_fpu_clock_0_out_waitrequest <= NOT nios2_fpu_clock_0_out_run;
  --nios2_fpu_clock_0_out_reset_n assignment, which is an e_assign
  nios2_fpu_clock_0_out_reset_n <= reset_n;
  --mux nios2_fpu_clock_0_out_endofpacket, which is an e_mux
  nios2_fpu_clock_0_out_endofpacket <= peripheral_bridge_s1_endofpacket_from_sa;
  --vhdl renameroo for output signals
  nios2_fpu_clock_0_out_address_to_slave <= internal_nios2_fpu_clock_0_out_address_to_slave;
  --vhdl renameroo for output signals
  nios2_fpu_clock_0_out_waitrequest <= internal_nios2_fpu_clock_0_out_waitrequest;
--synthesis translate_off
    --nios2_fpu_clock_0_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_clock_0_out_address_last_time <= std_logic_vector'("0000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_clock_0_out_address_last_time <= nios2_fpu_clock_0_out_address;
      end if;

    end process;

    --nios2_fpu_clock_0/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_nios2_fpu_clock_0_out_waitrequest AND ((nios2_fpu_clock_0_out_read OR nios2_fpu_clock_0_out_write));
      end if;

    end process;

    --nios2_fpu_clock_0_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line91 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_clock_0_out_address /= nios2_fpu_clock_0_out_address_last_time))))) = '1' then 
          write(write_line91, now);
          write(write_line91, string'(": "));
          write(write_line91, string'("nios2_fpu_clock_0_out_address did not heed wait!!!"));
          write(output, write_line91.all);
          deallocate (write_line91);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_clock_0_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_clock_0_out_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        nios2_fpu_clock_0_out_byteenable_last_time <= nios2_fpu_clock_0_out_byteenable;
      end if;

    end process;

    --nios2_fpu_clock_0_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line92 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_clock_0_out_byteenable /= nios2_fpu_clock_0_out_byteenable_last_time))))) = '1' then 
          write(write_line92, now);
          write(write_line92, string'(": "));
          write(write_line92, string'("nios2_fpu_clock_0_out_byteenable did not heed wait!!!"));
          write(output, write_line92.all);
          deallocate (write_line92);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_clock_0_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_clock_0_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_clock_0_out_read_last_time <= nios2_fpu_clock_0_out_read;
      end if;

    end process;

    --nios2_fpu_clock_0_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line93 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_clock_0_out_read) /= std_logic'(nios2_fpu_clock_0_out_read_last_time)))))) = '1' then 
          write(write_line93, now);
          write(write_line93, string'(": "));
          write(write_line93, string'("nios2_fpu_clock_0_out_read did not heed wait!!!"));
          write(output, write_line93.all);
          deallocate (write_line93);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_clock_0_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_clock_0_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        nios2_fpu_clock_0_out_write_last_time <= nios2_fpu_clock_0_out_write;
      end if;

    end process;

    --nios2_fpu_clock_0_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line94 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(nios2_fpu_clock_0_out_write) /= std_logic'(nios2_fpu_clock_0_out_write_last_time)))))) = '1' then 
          write(write_line94, now);
          write(write_line94, string'(": "));
          write(write_line94, string'("nios2_fpu_clock_0_out_write did not heed wait!!!"));
          write(output, write_line94.all);
          deallocate (write_line94);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_clock_0_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        nios2_fpu_clock_0_out_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        nios2_fpu_clock_0_out_writedata_last_time <= nios2_fpu_clock_0_out_writedata;
      end if;

    end process;

    --nios2_fpu_clock_0_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line95 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((nios2_fpu_clock_0_out_writedata /= nios2_fpu_clock_0_out_writedata_last_time)))) AND nios2_fpu_clock_0_out_write)) = '1' then 
          write(write_line95, now);
          write(write_line95, string'(": "));
          write(write_line95, string'("nios2_fpu_clock_0_out_writedata did not heed wait!!!"));
          write(output, write_line95.all);
          deallocate (write_line95);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_nios2_fpu_clock_0_out_to_peripheral_bridge_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_nios2_fpu_clock_0_out_to_peripheral_bridge_s1_module;


architecture europa of rdv_fifo_for_nios2_fpu_clock_0_out_to_peripheral_bridge_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (2 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_2;
  empty <= NOT(full_0);
  full_3 <= std_logic'('0');
  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 3);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 3);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 3);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity peripheral_bridge_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fpu_clock_0_out_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal nios2_fpu_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal nios2_fpu_clock_0_out_nativeaddress : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal nios2_fpu_clock_0_out_read : IN STD_LOGIC;
                 signal nios2_fpu_clock_0_out_write : IN STD_LOGIC;
                 signal nios2_fpu_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal peripheral_bridge_s1_endofpacket : IN STD_LOGIC;
                 signal peripheral_bridge_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal peripheral_bridge_s1_readdatavalid : IN STD_LOGIC;
                 signal peripheral_bridge_s1_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_peripheral_bridge_s1_end_xfer : OUT STD_LOGIC;
                 signal nios2_fpu_clock_0_out_granted_peripheral_bridge_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1_shift_register : OUT STD_LOGIC;
                 signal nios2_fpu_clock_0_out_requests_peripheral_bridge_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_s1_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal peripheral_bridge_s1_arbiterlock : OUT STD_LOGIC;
                 signal peripheral_bridge_s1_arbiterlock2 : OUT STD_LOGIC;
                 signal peripheral_bridge_s1_burstcount : OUT STD_LOGIC;
                 signal peripheral_bridge_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal peripheral_bridge_s1_chipselect : OUT STD_LOGIC;
                 signal peripheral_bridge_s1_debugaccess : OUT STD_LOGIC;
                 signal peripheral_bridge_s1_endofpacket_from_sa : OUT STD_LOGIC;
                 signal peripheral_bridge_s1_nativeaddress : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal peripheral_bridge_s1_read : OUT STD_LOGIC;
                 signal peripheral_bridge_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal peripheral_bridge_s1_reset_n : OUT STD_LOGIC;
                 signal peripheral_bridge_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal peripheral_bridge_s1_write : OUT STD_LOGIC;
                 signal peripheral_bridge_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity peripheral_bridge_s1_arbitrator;


architecture europa of peripheral_bridge_s1_arbitrator is
component rdv_fifo_for_nios2_fpu_clock_0_out_to_peripheral_bridge_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_nios2_fpu_clock_0_out_to_peripheral_bridge_s1_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_peripheral_bridge_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_fpu_clock_0_out_granted_peripheral_bridge_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1_shift_register :  STD_LOGIC;
                signal internal_nios2_fpu_clock_0_out_requests_peripheral_bridge_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_s1_waitrequest_from_sa :  STD_LOGIC;
                signal module_input54 :  STD_LOGIC;
                signal module_input55 :  STD_LOGIC;
                signal module_input56 :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_arbiterlock :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_arbiterlock2 :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_continuerequest :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_rdv_fifo_empty_peripheral_bridge_s1 :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_rdv_fifo_output_from_peripheral_bridge_s1 :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_saved_grant_peripheral_bridge_s1 :  STD_LOGIC;
                signal peripheral_bridge_s1_allgrants :  STD_LOGIC;
                signal peripheral_bridge_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal peripheral_bridge_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal peripheral_bridge_s1_any_continuerequest :  STD_LOGIC;
                signal peripheral_bridge_s1_arb_counter_enable :  STD_LOGIC;
                signal peripheral_bridge_s1_arb_share_counter :  STD_LOGIC;
                signal peripheral_bridge_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal peripheral_bridge_s1_arb_share_set_values :  STD_LOGIC;
                signal peripheral_bridge_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal peripheral_bridge_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal peripheral_bridge_s1_begins_xfer :  STD_LOGIC;
                signal peripheral_bridge_s1_end_xfer :  STD_LOGIC;
                signal peripheral_bridge_s1_firsttransfer :  STD_LOGIC;
                signal peripheral_bridge_s1_grant_vector :  STD_LOGIC;
                signal peripheral_bridge_s1_in_a_read_cycle :  STD_LOGIC;
                signal peripheral_bridge_s1_in_a_write_cycle :  STD_LOGIC;
                signal peripheral_bridge_s1_master_qreq_vector :  STD_LOGIC;
                signal peripheral_bridge_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal peripheral_bridge_s1_non_bursting_master_requests :  STD_LOGIC;
                signal peripheral_bridge_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal peripheral_bridge_s1_reg_firsttransfer :  STD_LOGIC;
                signal peripheral_bridge_s1_slavearbiterlockenable :  STD_LOGIC;
                signal peripheral_bridge_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal peripheral_bridge_s1_unreg_firsttransfer :  STD_LOGIC;
                signal peripheral_bridge_s1_waits_for_read :  STD_LOGIC;
                signal peripheral_bridge_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_peripheral_bridge_s1_from_nios2_fpu_clock_0_out :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal wait_for_peripheral_bridge_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT peripheral_bridge_s1_end_xfer;
    end if;

  end process;

  peripheral_bridge_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1);
  --assign peripheral_bridge_s1_readdata_from_sa = peripheral_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  peripheral_bridge_s1_readdata_from_sa <= peripheral_bridge_s1_readdata;
  internal_nios2_fpu_clock_0_out_requests_peripheral_bridge_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_clock_0_out_read OR nios2_fpu_clock_0_out_write)))))));
  --assign peripheral_bridge_s1_waitrequest_from_sa = peripheral_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_peripheral_bridge_s1_waitrequest_from_sa <= peripheral_bridge_s1_waitrequest;
  --assign peripheral_bridge_s1_readdatavalid_from_sa = peripheral_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  peripheral_bridge_s1_readdatavalid_from_sa <= peripheral_bridge_s1_readdatavalid;
  --peripheral_bridge_s1_arb_share_counter set values, which is an e_mux
  peripheral_bridge_s1_arb_share_set_values <= std_logic'('1');
  --peripheral_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  peripheral_bridge_s1_non_bursting_master_requests <= internal_nios2_fpu_clock_0_out_requests_peripheral_bridge_s1 OR internal_nios2_fpu_clock_0_out_requests_peripheral_bridge_s1;
  --peripheral_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  peripheral_bridge_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --peripheral_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  peripheral_bridge_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(peripheral_bridge_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(peripheral_bridge_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --peripheral_bridge_s1_allgrants all slave grants, which is an e_mux
  peripheral_bridge_s1_allgrants <= (peripheral_bridge_s1_grant_vector) OR (peripheral_bridge_s1_grant_vector);
  --peripheral_bridge_s1_end_xfer assignment, which is an e_assign
  peripheral_bridge_s1_end_xfer <= NOT ((peripheral_bridge_s1_waits_for_read OR peripheral_bridge_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_peripheral_bridge_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_peripheral_bridge_s1 <= peripheral_bridge_s1_end_xfer AND (((NOT peripheral_bridge_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --peripheral_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  peripheral_bridge_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_peripheral_bridge_s1 AND peripheral_bridge_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_peripheral_bridge_s1 AND NOT peripheral_bridge_s1_non_bursting_master_requests));
  --peripheral_bridge_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      peripheral_bridge_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(peripheral_bridge_s1_arb_counter_enable) = '1' then 
        peripheral_bridge_s1_arb_share_counter <= peripheral_bridge_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --peripheral_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      peripheral_bridge_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((peripheral_bridge_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_peripheral_bridge_s1)) OR ((end_xfer_arb_share_counter_term_peripheral_bridge_s1 AND NOT peripheral_bridge_s1_non_bursting_master_requests)))) = '1' then 
        peripheral_bridge_s1_slavearbiterlockenable <= peripheral_bridge_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --nios2_fpu_clock_0/out peripheral_bridge/s1 arbiterlock, which is an e_assign
  nios2_fpu_clock_0_out_arbiterlock <= peripheral_bridge_s1_slavearbiterlockenable AND nios2_fpu_clock_0_out_continuerequest;
  --peripheral_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  peripheral_bridge_s1_slavearbiterlockenable2 <= peripheral_bridge_s1_arb_share_counter_next_value;
  --nios2_fpu_clock_0/out peripheral_bridge/s1 arbiterlock2, which is an e_assign
  nios2_fpu_clock_0_out_arbiterlock2 <= peripheral_bridge_s1_slavearbiterlockenable2 AND nios2_fpu_clock_0_out_continuerequest;
  --peripheral_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  peripheral_bridge_s1_any_continuerequest <= std_logic'('1');
  --nios2_fpu_clock_0_out_continuerequest continued request, which is an e_assign
  nios2_fpu_clock_0_out_continuerequest <= std_logic'('1');
  internal_nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1 <= internal_nios2_fpu_clock_0_out_requests_peripheral_bridge_s1 AND NOT ((nios2_fpu_clock_0_out_read AND (internal_nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1_shift_register)));
  --unique name for peripheral_bridge_s1_move_on_to_next_transaction, which is an e_assign
  peripheral_bridge_s1_move_on_to_next_transaction <= peripheral_bridge_s1_readdatavalid_from_sa;
  --rdv_fifo_for_nios2_fpu_clock_0_out_to_peripheral_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios2_fpu_clock_0_out_to_peripheral_bridge_s1 : rdv_fifo_for_nios2_fpu_clock_0_out_to_peripheral_bridge_s1_module
    port map(
      data_out => nios2_fpu_clock_0_out_rdv_fifo_output_from_peripheral_bridge_s1,
      empty => open,
      fifo_contains_ones_n => nios2_fpu_clock_0_out_rdv_fifo_empty_peripheral_bridge_s1,
      full => open,
      clear_fifo => module_input54,
      clk => clk,
      data_in => internal_nios2_fpu_clock_0_out_granted_peripheral_bridge_s1,
      read => peripheral_bridge_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input55,
      write => module_input56
    );

  module_input54 <= std_logic'('0');
  module_input55 <= std_logic'('0');
  module_input56 <= in_a_read_cycle AND NOT peripheral_bridge_s1_waits_for_read;

  internal_nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1_shift_register <= NOT nios2_fpu_clock_0_out_rdv_fifo_empty_peripheral_bridge_s1;
  --local readdatavalid nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1, which is an e_mux
  nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1 <= peripheral_bridge_s1_readdatavalid_from_sa;
  --peripheral_bridge_s1_writedata mux, which is an e_mux
  peripheral_bridge_s1_writedata <= nios2_fpu_clock_0_out_writedata;
  --assign peripheral_bridge_s1_endofpacket_from_sa = peripheral_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  peripheral_bridge_s1_endofpacket_from_sa <= peripheral_bridge_s1_endofpacket;
  --master is always granted when requested
  internal_nios2_fpu_clock_0_out_granted_peripheral_bridge_s1 <= internal_nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1;
  --nios2_fpu_clock_0/out saved-grant peripheral_bridge/s1, which is an e_assign
  nios2_fpu_clock_0_out_saved_grant_peripheral_bridge_s1 <= internal_nios2_fpu_clock_0_out_requests_peripheral_bridge_s1;
  --allow new arb cycle for peripheral_bridge/s1, which is an e_assign
  peripheral_bridge_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  peripheral_bridge_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  peripheral_bridge_s1_master_qreq_vector <= std_logic'('1');
  --peripheral_bridge_s1_reset_n assignment, which is an e_assign
  peripheral_bridge_s1_reset_n <= reset_n;
  peripheral_bridge_s1_chipselect <= internal_nios2_fpu_clock_0_out_granted_peripheral_bridge_s1;
  --peripheral_bridge_s1_firsttransfer first transaction, which is an e_assign
  peripheral_bridge_s1_firsttransfer <= A_WE_StdLogic((std_logic'(peripheral_bridge_s1_begins_xfer) = '1'), peripheral_bridge_s1_unreg_firsttransfer, peripheral_bridge_s1_reg_firsttransfer);
  --peripheral_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  peripheral_bridge_s1_unreg_firsttransfer <= NOT ((peripheral_bridge_s1_slavearbiterlockenable AND peripheral_bridge_s1_any_continuerequest));
  --peripheral_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      peripheral_bridge_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(peripheral_bridge_s1_begins_xfer) = '1' then 
        peripheral_bridge_s1_reg_firsttransfer <= peripheral_bridge_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --peripheral_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  peripheral_bridge_s1_beginbursttransfer_internal <= peripheral_bridge_s1_begins_xfer;
  --peripheral_bridge_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  peripheral_bridge_s1_arbitration_holdoff_internal <= peripheral_bridge_s1_begins_xfer AND peripheral_bridge_s1_firsttransfer;
  --peripheral_bridge_s1_read assignment, which is an e_mux
  peripheral_bridge_s1_read <= internal_nios2_fpu_clock_0_out_granted_peripheral_bridge_s1 AND nios2_fpu_clock_0_out_read;
  --peripheral_bridge_s1_write assignment, which is an e_mux
  peripheral_bridge_s1_write <= internal_nios2_fpu_clock_0_out_granted_peripheral_bridge_s1 AND nios2_fpu_clock_0_out_write;
  shifted_address_to_peripheral_bridge_s1_from_nios2_fpu_clock_0_out <= nios2_fpu_clock_0_out_address_to_slave;
  --peripheral_bridge_s1_address mux, which is an e_mux
  peripheral_bridge_s1_address <= A_EXT (A_SRL(shifted_address_to_peripheral_bridge_s1_from_nios2_fpu_clock_0_out,std_logic_vector'("00000000000000000000000000000010")), 11);
  --slaveid peripheral_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  peripheral_bridge_s1_nativeaddress <= nios2_fpu_clock_0_out_nativeaddress;
  --d1_peripheral_bridge_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_peripheral_bridge_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_peripheral_bridge_s1_end_xfer <= peripheral_bridge_s1_end_xfer;
    end if;

  end process;

  --peripheral_bridge_s1_waits_for_read in a cycle, which is an e_mux
  peripheral_bridge_s1_waits_for_read <= peripheral_bridge_s1_in_a_read_cycle AND internal_peripheral_bridge_s1_waitrequest_from_sa;
  --peripheral_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  peripheral_bridge_s1_in_a_read_cycle <= internal_nios2_fpu_clock_0_out_granted_peripheral_bridge_s1 AND nios2_fpu_clock_0_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= peripheral_bridge_s1_in_a_read_cycle;
  --peripheral_bridge_s1_waits_for_write in a cycle, which is an e_mux
  peripheral_bridge_s1_waits_for_write <= peripheral_bridge_s1_in_a_write_cycle AND internal_peripheral_bridge_s1_waitrequest_from_sa;
  --peripheral_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  peripheral_bridge_s1_in_a_write_cycle <= internal_nios2_fpu_clock_0_out_granted_peripheral_bridge_s1 AND nios2_fpu_clock_0_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= peripheral_bridge_s1_in_a_write_cycle;
  wait_for_peripheral_bridge_s1_counter <= std_logic'('0');
  --peripheral_bridge_s1_byteenable byte enable port mux, which is an e_mux
  peripheral_bridge_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_clock_0_out_granted_peripheral_bridge_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (nios2_fpu_clock_0_out_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --burstcount mux, which is an e_mux
  peripheral_bridge_s1_burstcount <= std_logic'('1');
  --peripheral_bridge/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  peripheral_bridge_s1_arbiterlock <= nios2_fpu_clock_0_out_arbiterlock;
  --peripheral_bridge/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  peripheral_bridge_s1_arbiterlock2 <= nios2_fpu_clock_0_out_arbiterlock2;
  --debugaccess mux, which is an e_mux
  peripheral_bridge_s1_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  nios2_fpu_clock_0_out_granted_peripheral_bridge_s1 <= internal_nios2_fpu_clock_0_out_granted_peripheral_bridge_s1;
  --vhdl renameroo for output signals
  nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1 <= internal_nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1;
  --vhdl renameroo for output signals
  nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1_shift_register <= internal_nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1_shift_register;
  --vhdl renameroo for output signals
  nios2_fpu_clock_0_out_requests_peripheral_bridge_s1 <= internal_nios2_fpu_clock_0_out_requests_peripheral_bridge_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_s1_waitrequest_from_sa <= internal_peripheral_bridge_s1_waitrequest_from_sa;
--synthesis translate_off
    --peripheral_bridge/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity peripheral_bridge_m1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_dipsw_s1_end_xfer : IN STD_LOGIC;
                 signal d1_gpio0_s1_end_xfer : IN STD_LOGIC;
                 signal d1_jtag_uart_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                 signal d1_led_s1_end_xfer : IN STD_LOGIC;
                 signal d1_mmcdma_s1_end_xfer : IN STD_LOGIC;
                 signal d1_psw_s1_end_xfer : IN STD_LOGIC;
                 signal d1_spu_s1_end_xfer : IN STD_LOGIC;
                 signal d1_sysid_control_slave_end_xfer : IN STD_LOGIC;
                 signal d1_systimer_s1_end_xfer : IN STD_LOGIC;
                 signal d1_sysuart_s1_end_xfer : IN STD_LOGIC;
                 signal d1_vga_s1_end_xfer : IN STD_LOGIC;
                 signal dipsw_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal gpio0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal led_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal mmcdma_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal mmcdma_s1_wait_counter_eq_0 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                 signal peripheral_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                 signal peripheral_bridge_m1_granted_dipsw_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_granted_gpio0_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal peripheral_bridge_m1_granted_led_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_granted_mmcdma_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_granted_psw_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_granted_spu_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_granted_sysid_control_slave : IN STD_LOGIC;
                 signal peripheral_bridge_m1_granted_systimer_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_granted_sysuart_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_granted_vga_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_dipsw_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_gpio0_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_led_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_mmcdma_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_psw_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_spu_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_sysid_control_slave : IN STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_systimer_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_sysuart_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_vga_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_dipsw_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_gpio0_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_led_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_mmcdma_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_psw_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_spu_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_sysid_control_slave : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_systimer_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_sysuart_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_vga_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_requests_dipsw_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_requests_gpio0_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal peripheral_bridge_m1_requests_led_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_requests_mmcdma_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_requests_psw_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_requests_spu_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_requests_sysid_control_slave : IN STD_LOGIC;
                 signal peripheral_bridge_m1_requests_systimer_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_requests_sysuart_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_requests_vga_s1 : IN STD_LOGIC;
                 signal peripheral_bridge_m1_write : IN STD_LOGIC;
                 signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal psw_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal spu_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal spu_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal sysid_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal systimer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sysuart_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal vga_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal peripheral_bridge_m1_address_to_slave : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal peripheral_bridge_m1_latency_counter : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal peripheral_bridge_m1_readdatavalid : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_waitrequest : OUT STD_LOGIC
              );
end entity peripheral_bridge_m1_arbitrator;


architecture europa of peripheral_bridge_m1_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_address_to_slave :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal internal_peripheral_bridge_m1_latency_counter :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal p1_peripheral_bridge_m1_latency_counter :  STD_LOGIC;
                signal peripheral_bridge_m1_address_last_time :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal peripheral_bridge_m1_burstcount_last_time :  STD_LOGIC;
                signal peripheral_bridge_m1_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal peripheral_bridge_m1_chipselect_last_time :  STD_LOGIC;
                signal peripheral_bridge_m1_is_granted_some_slave :  STD_LOGIC;
                signal peripheral_bridge_m1_read_but_no_slave_selected :  STD_LOGIC;
                signal peripheral_bridge_m1_read_last_time :  STD_LOGIC;
                signal peripheral_bridge_m1_run :  STD_LOGIC;
                signal peripheral_bridge_m1_write_last_time :  STD_LOGIC;
                signal peripheral_bridge_m1_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pre_flush_peripheral_bridge_m1_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_qualified_request_dipsw_s1 OR NOT peripheral_bridge_m1_requests_dipsw_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_dipsw_s1 OR NOT ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_dipsw_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_dipsw_s1 OR NOT ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_qualified_request_gpio0_s1 OR NOT peripheral_bridge_m1_requests_gpio0_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_gpio0_s1 OR NOT ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_gpio0_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_gpio0_s1 OR NOT ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave OR NOT peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave OR NOT peripheral_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_chipselect)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave OR NOT peripheral_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_chipselect)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_qualified_request_led_s1 OR NOT peripheral_bridge_m1_requests_led_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_led_s1 OR NOT ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_led_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_led_s1 OR NOT ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_qualified_request_mmcdma_s1 OR NOT peripheral_bridge_m1_requests_mmcdma_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_mmcdma_s1 OR NOT ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((mmcdma_s1_wait_counter_eq_0 AND NOT d1_mmcdma_s1_end_xfer)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_mmcdma_s1 OR NOT ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))))))));
  --cascaded wait assignment, which is an e_assign
  peripheral_bridge_m1_run <= (r_0 AND r_1) AND r_2;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_qualified_request_psw_s1 OR NOT peripheral_bridge_m1_requests_psw_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_psw_s1 OR NOT ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_psw_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_psw_s1 OR NOT ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_qualified_request_spu_s1 OR NOT peripheral_bridge_m1_requests_spu_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_spu_s1 OR NOT peripheral_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT spu_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_chipselect)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_spu_s1 OR NOT peripheral_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT spu_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_chipselect)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_qualified_request_sysid_control_slave OR NOT peripheral_bridge_m1_requests_sysid_control_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_sysid_control_slave OR NOT ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_sysid_control_slave_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_sysid_control_slave OR NOT ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_qualified_request_systimer_s1 OR NOT peripheral_bridge_m1_requests_systimer_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_systimer_s1 OR NOT ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_systimer_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_systimer_s1 OR NOT ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_qualified_request_sysuart_s1 OR NOT peripheral_bridge_m1_requests_sysuart_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_sysuart_s1 OR NOT peripheral_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_sysuart_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_chipselect)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_sysuart_s1 OR NOT peripheral_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_sysuart_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_chipselect)))))))));
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_qualified_request_vga_s1 OR NOT peripheral_bridge_m1_requests_vga_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_vga_s1 OR NOT ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_vga_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT peripheral_bridge_m1_qualified_request_vga_s1 OR NOT ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_peripheral_bridge_m1_address_to_slave <= peripheral_bridge_m1_address(12 DOWNTO 0);
  --peripheral_bridge_m1_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      peripheral_bridge_m1_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      peripheral_bridge_m1_read_but_no_slave_selected <= (((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)) AND peripheral_bridge_m1_run) AND NOT peripheral_bridge_m1_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  peripheral_bridge_m1_is_granted_some_slave <= (((((((((peripheral_bridge_m1_granted_dipsw_s1 OR peripheral_bridge_m1_granted_gpio0_s1) OR peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave) OR peripheral_bridge_m1_granted_led_s1) OR peripheral_bridge_m1_granted_mmcdma_s1) OR peripheral_bridge_m1_granted_psw_s1) OR peripheral_bridge_m1_granted_spu_s1) OR peripheral_bridge_m1_granted_sysid_control_slave) OR peripheral_bridge_m1_granted_systimer_s1) OR peripheral_bridge_m1_granted_sysuart_s1) OR peripheral_bridge_m1_granted_vga_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_peripheral_bridge_m1_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  peripheral_bridge_m1_readdatavalid <= (((((((((((((((((((((((((((((((peripheral_bridge_m1_read_but_no_slave_selected OR pre_flush_peripheral_bridge_m1_readdatavalid) OR peripheral_bridge_m1_read_data_valid_dipsw_s1) OR peripheral_bridge_m1_read_but_no_slave_selected) OR pre_flush_peripheral_bridge_m1_readdatavalid) OR peripheral_bridge_m1_read_data_valid_gpio0_s1) OR peripheral_bridge_m1_read_but_no_slave_selected) OR pre_flush_peripheral_bridge_m1_readdatavalid) OR peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave) OR peripheral_bridge_m1_read_but_no_slave_selected) OR pre_flush_peripheral_bridge_m1_readdatavalid) OR peripheral_bridge_m1_read_data_valid_led_s1) OR peripheral_bridge_m1_read_but_no_slave_selected) OR pre_flush_peripheral_bridge_m1_readdatavalid) OR peripheral_bridge_m1_read_data_valid_mmcdma_s1) OR peripheral_bridge_m1_read_but_no_slave_selected) OR pre_flush_peripheral_bridge_m1_readdatavalid) OR peripheral_bridge_m1_read_data_valid_psw_s1) OR peripheral_bridge_m1_read_but_no_slave_selected) OR pre_flush_peripheral_bridge_m1_readdatavalid) OR peripheral_bridge_m1_read_data_valid_spu_s1) OR peripheral_bridge_m1_read_but_no_slave_selected) OR pre_flush_peripheral_bridge_m1_readdatavalid) OR peripheral_bridge_m1_read_data_valid_sysid_control_slave) OR peripheral_bridge_m1_read_but_no_slave_selected) OR pre_flush_peripheral_bridge_m1_readdatavalid) OR peripheral_bridge_m1_read_data_valid_systimer_s1) OR peripheral_bridge_m1_read_but_no_slave_selected) OR pre_flush_peripheral_bridge_m1_readdatavalid) OR peripheral_bridge_m1_read_data_valid_sysuart_s1) OR peripheral_bridge_m1_read_but_no_slave_selected) OR pre_flush_peripheral_bridge_m1_readdatavalid) OR peripheral_bridge_m1_read_data_valid_vga_s1;
  --peripheral_bridge/m1 readdata mux, which is an e_mux
  peripheral_bridge_m1_readdata <= (((((((((((A_REP(NOT ((peripheral_bridge_m1_qualified_request_dipsw_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))) , 32) OR dipsw_s1_readdata_from_sa)) AND ((A_REP(NOT ((peripheral_bridge_m1_qualified_request_gpio0_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))) , 32) OR gpio0_s1_readdata_from_sa))) AND ((A_REP(NOT ((peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))) , 32) OR jtag_uart_avalon_jtag_slave_readdata_from_sa))) AND ((A_REP(NOT ((peripheral_bridge_m1_qualified_request_led_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))) , 32) OR led_s1_readdata_from_sa))) AND ((A_REP(NOT ((peripheral_bridge_m1_qualified_request_mmcdma_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))) , 32) OR mmcdma_s1_readdata_from_sa))) AND ((A_REP(NOT ((peripheral_bridge_m1_qualified_request_psw_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))) , 32) OR psw_s1_readdata_from_sa))) AND ((A_REP(NOT ((peripheral_bridge_m1_qualified_request_spu_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))) , 32) OR spu_s1_readdata_from_sa))) AND ((A_REP(NOT ((peripheral_bridge_m1_qualified_request_sysid_control_slave AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))) , 32) OR sysid_control_slave_readdata_from_sa))) AND ((A_REP(NOT ((peripheral_bridge_m1_qualified_request_systimer_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))) , 32) OR (std_logic_vector'("0000000000000000") & (systimer_s1_readdata_from_sa))))) AND ((A_REP(NOT ((peripheral_bridge_m1_qualified_request_sysuart_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))) , 32) OR (std_logic_vector'("0000000000000000") & (sysuart_s1_readdata_from_sa))))) AND ((A_REP(NOT ((peripheral_bridge_m1_qualified_request_vga_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)))) , 32) OR vga_s1_readdata_from_sa));
  --actual waitrequest port, which is an e_assign
  internal_peripheral_bridge_m1_waitrequest <= NOT peripheral_bridge_m1_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_peripheral_bridge_m1_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_peripheral_bridge_m1_latency_counter <= p1_peripheral_bridge_m1_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_peripheral_bridge_m1_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((peripheral_bridge_m1_run AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect))))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_peripheral_bridge_m1_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_peripheral_bridge_m1_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --vhdl renameroo for output signals
  peripheral_bridge_m1_address_to_slave <= internal_peripheral_bridge_m1_address_to_slave;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_latency_counter <= internal_peripheral_bridge_m1_latency_counter;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_waitrequest <= internal_peripheral_bridge_m1_waitrequest;
--synthesis translate_off
    --peripheral_bridge_m1_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        peripheral_bridge_m1_address_last_time <= std_logic_vector'("0000000000000");
      elsif clk'event and clk = '1' then
        peripheral_bridge_m1_address_last_time <= peripheral_bridge_m1_address;
      end if;

    end process;

    --peripheral_bridge/m1 waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_peripheral_bridge_m1_waitrequest AND peripheral_bridge_m1_chipselect;
      end if;

    end process;

    --peripheral_bridge_m1_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line96 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((peripheral_bridge_m1_address /= peripheral_bridge_m1_address_last_time))))) = '1' then 
          write(write_line96, now);
          write(write_line96, string'(": "));
          write(write_line96, string'("peripheral_bridge_m1_address did not heed wait!!!"));
          write(output, write_line96.all);
          deallocate (write_line96);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --peripheral_bridge_m1_chipselect check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        peripheral_bridge_m1_chipselect_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        peripheral_bridge_m1_chipselect_last_time <= peripheral_bridge_m1_chipselect;
      end if;

    end process;

    --peripheral_bridge_m1_chipselect matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line97 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(peripheral_bridge_m1_chipselect) /= std_logic'(peripheral_bridge_m1_chipselect_last_time)))))) = '1' then 
          write(write_line97, now);
          write(write_line97, string'(": "));
          write(write_line97, string'("peripheral_bridge_m1_chipselect did not heed wait!!!"));
          write(output, write_line97.all);
          deallocate (write_line97);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --peripheral_bridge_m1_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        peripheral_bridge_m1_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        peripheral_bridge_m1_burstcount_last_time <= peripheral_bridge_m1_burstcount;
      end if;

    end process;

    --peripheral_bridge_m1_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line98 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(peripheral_bridge_m1_burstcount) /= std_logic'(peripheral_bridge_m1_burstcount_last_time)))))) = '1' then 
          write(write_line98, now);
          write(write_line98, string'(": "));
          write(write_line98, string'("peripheral_bridge_m1_burstcount did not heed wait!!!"));
          write(output, write_line98.all);
          deallocate (write_line98);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --peripheral_bridge_m1_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        peripheral_bridge_m1_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        peripheral_bridge_m1_byteenable_last_time <= peripheral_bridge_m1_byteenable;
      end if;

    end process;

    --peripheral_bridge_m1_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line99 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((peripheral_bridge_m1_byteenable /= peripheral_bridge_m1_byteenable_last_time))))) = '1' then 
          write(write_line99, now);
          write(write_line99, string'(": "));
          write(write_line99, string'("peripheral_bridge_m1_byteenable did not heed wait!!!"));
          write(output, write_line99.all);
          deallocate (write_line99);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --peripheral_bridge_m1_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        peripheral_bridge_m1_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        peripheral_bridge_m1_read_last_time <= peripheral_bridge_m1_read;
      end if;

    end process;

    --peripheral_bridge_m1_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line100 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(peripheral_bridge_m1_read) /= std_logic'(peripheral_bridge_m1_read_last_time)))))) = '1' then 
          write(write_line100, now);
          write(write_line100, string'(": "));
          write(write_line100, string'("peripheral_bridge_m1_read did not heed wait!!!"));
          write(output, write_line100.all);
          deallocate (write_line100);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --peripheral_bridge_m1_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        peripheral_bridge_m1_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        peripheral_bridge_m1_write_last_time <= peripheral_bridge_m1_write;
      end if;

    end process;

    --peripheral_bridge_m1_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line101 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(peripheral_bridge_m1_write) /= std_logic'(peripheral_bridge_m1_write_last_time)))))) = '1' then 
          write(write_line101, now);
          write(write_line101, string'(": "));
          write(write_line101, string'("peripheral_bridge_m1_write did not heed wait!!!"));
          write(output, write_line101.all);
          deallocate (write_line101);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --peripheral_bridge_m1_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        peripheral_bridge_m1_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        peripheral_bridge_m1_writedata_last_time <= peripheral_bridge_m1_writedata;
      end if;

    end process;

    --peripheral_bridge_m1_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line102 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((peripheral_bridge_m1_writedata /= peripheral_bridge_m1_writedata_last_time)))) AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect)))) = '1' then 
          write(write_line102, now);
          write(write_line102, string'(": "));
          write(write_line102, string'("peripheral_bridge_m1_writedata did not heed wait!!!"));
          write(output, write_line102.all);
          deallocate (write_line102);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity peripheral_bridge_bridge_arbitrator is 
end entity peripheral_bridge_bridge_arbitrator;


architecture europa of peripheral_bridge_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity psw_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                 signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                 signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read : IN STD_LOGIC;
                 signal peripheral_bridge_m1_write : IN STD_LOGIC;
                 signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal psw_s1_irq : IN STD_LOGIC;
                 signal psw_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_psw_s1_end_xfer : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_granted_psw_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_psw_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_psw_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_requests_psw_s1 : OUT STD_LOGIC;
                 signal psw_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal psw_s1_chipselect : OUT STD_LOGIC;
                 signal psw_s1_irq_from_sa : OUT STD_LOGIC;
                 signal psw_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal psw_s1_reset_n : OUT STD_LOGIC;
                 signal psw_s1_write_n : OUT STD_LOGIC;
                 signal psw_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity psw_s1_arbitrator;


architecture europa of psw_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_psw_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_granted_psw_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_qualified_request_psw_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_requests_psw_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal peripheral_bridge_m1_continuerequest :  STD_LOGIC;
                signal peripheral_bridge_m1_saved_grant_psw_s1 :  STD_LOGIC;
                signal psw_s1_allgrants :  STD_LOGIC;
                signal psw_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal psw_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal psw_s1_any_continuerequest :  STD_LOGIC;
                signal psw_s1_arb_counter_enable :  STD_LOGIC;
                signal psw_s1_arb_share_counter :  STD_LOGIC;
                signal psw_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal psw_s1_arb_share_set_values :  STD_LOGIC;
                signal psw_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal psw_s1_begins_xfer :  STD_LOGIC;
                signal psw_s1_end_xfer :  STD_LOGIC;
                signal psw_s1_firsttransfer :  STD_LOGIC;
                signal psw_s1_grant_vector :  STD_LOGIC;
                signal psw_s1_in_a_read_cycle :  STD_LOGIC;
                signal psw_s1_in_a_write_cycle :  STD_LOGIC;
                signal psw_s1_master_qreq_vector :  STD_LOGIC;
                signal psw_s1_non_bursting_master_requests :  STD_LOGIC;
                signal psw_s1_reg_firsttransfer :  STD_LOGIC;
                signal psw_s1_slavearbiterlockenable :  STD_LOGIC;
                signal psw_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal psw_s1_unreg_firsttransfer :  STD_LOGIC;
                signal psw_s1_waits_for_read :  STD_LOGIC;
                signal psw_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_psw_s1_from_peripheral_bridge_m1 :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal wait_for_psw_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT psw_s1_end_xfer;
    end if;

  end process;

  psw_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_peripheral_bridge_m1_qualified_request_psw_s1);
  --assign psw_s1_readdata_from_sa = psw_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  psw_s1_readdata_from_sa <= psw_s1_readdata;
  internal_peripheral_bridge_m1_requests_psw_s1 <= to_std_logic(((Std_Logic_Vector'(peripheral_bridge_m1_address_to_slave(12 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("0001001000000")))) AND peripheral_bridge_m1_chipselect;
  --psw_s1_arb_share_counter set values, which is an e_mux
  psw_s1_arb_share_set_values <= std_logic'('1');
  --psw_s1_non_bursting_master_requests mux, which is an e_mux
  psw_s1_non_bursting_master_requests <= internal_peripheral_bridge_m1_requests_psw_s1;
  --psw_s1_any_bursting_master_saved_grant mux, which is an e_mux
  psw_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --psw_s1_arb_share_counter_next_value assignment, which is an e_assign
  psw_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(psw_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(psw_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(psw_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(psw_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --psw_s1_allgrants all slave grants, which is an e_mux
  psw_s1_allgrants <= psw_s1_grant_vector;
  --psw_s1_end_xfer assignment, which is an e_assign
  psw_s1_end_xfer <= NOT ((psw_s1_waits_for_read OR psw_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_psw_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_psw_s1 <= psw_s1_end_xfer AND (((NOT psw_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --psw_s1_arb_share_counter arbitration counter enable, which is an e_assign
  psw_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_psw_s1 AND psw_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_psw_s1 AND NOT psw_s1_non_bursting_master_requests));
  --psw_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      psw_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(psw_s1_arb_counter_enable) = '1' then 
        psw_s1_arb_share_counter <= psw_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --psw_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      psw_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((psw_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_psw_s1)) OR ((end_xfer_arb_share_counter_term_psw_s1 AND NOT psw_s1_non_bursting_master_requests)))) = '1' then 
        psw_s1_slavearbiterlockenable <= psw_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --peripheral_bridge/m1 psw/s1 arbiterlock, which is an e_assign
  peripheral_bridge_m1_arbiterlock <= psw_s1_slavearbiterlockenable AND peripheral_bridge_m1_continuerequest;
  --psw_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  psw_s1_slavearbiterlockenable2 <= psw_s1_arb_share_counter_next_value;
  --peripheral_bridge/m1 psw/s1 arbiterlock2, which is an e_assign
  peripheral_bridge_m1_arbiterlock2 <= psw_s1_slavearbiterlockenable2 AND peripheral_bridge_m1_continuerequest;
  --psw_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  psw_s1_any_continuerequest <= std_logic'('1');
  --peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  peripheral_bridge_m1_continuerequest <= std_logic'('1');
  internal_peripheral_bridge_m1_qualified_request_psw_s1 <= internal_peripheral_bridge_m1_requests_psw_s1 AND NOT ((((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid peripheral_bridge_m1_read_data_valid_psw_s1, which is an e_mux
  peripheral_bridge_m1_read_data_valid_psw_s1 <= (internal_peripheral_bridge_m1_granted_psw_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect))) AND NOT psw_s1_waits_for_read;
  --psw_s1_writedata mux, which is an e_mux
  psw_s1_writedata <= peripheral_bridge_m1_writedata;
  --master is always granted when requested
  internal_peripheral_bridge_m1_granted_psw_s1 <= internal_peripheral_bridge_m1_qualified_request_psw_s1;
  --peripheral_bridge/m1 saved-grant psw/s1, which is an e_assign
  peripheral_bridge_m1_saved_grant_psw_s1 <= internal_peripheral_bridge_m1_requests_psw_s1;
  --allow new arb cycle for psw/s1, which is an e_assign
  psw_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  psw_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  psw_s1_master_qreq_vector <= std_logic'('1');
  --psw_s1_reset_n assignment, which is an e_assign
  psw_s1_reset_n <= reset_n;
  psw_s1_chipselect <= internal_peripheral_bridge_m1_granted_psw_s1;
  --psw_s1_firsttransfer first transaction, which is an e_assign
  psw_s1_firsttransfer <= A_WE_StdLogic((std_logic'(psw_s1_begins_xfer) = '1'), psw_s1_unreg_firsttransfer, psw_s1_reg_firsttransfer);
  --psw_s1_unreg_firsttransfer first transaction, which is an e_assign
  psw_s1_unreg_firsttransfer <= NOT ((psw_s1_slavearbiterlockenable AND psw_s1_any_continuerequest));
  --psw_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      psw_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(psw_s1_begins_xfer) = '1' then 
        psw_s1_reg_firsttransfer <= psw_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --psw_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  psw_s1_beginbursttransfer_internal <= psw_s1_begins_xfer;
  --~psw_s1_write_n assignment, which is an e_mux
  psw_s1_write_n <= NOT ((internal_peripheral_bridge_m1_granted_psw_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect))));
  shifted_address_to_psw_s1_from_peripheral_bridge_m1 <= peripheral_bridge_m1_address_to_slave;
  --psw_s1_address mux, which is an e_mux
  psw_s1_address <= A_EXT (A_SRL(shifted_address_to_psw_s1_from_peripheral_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_psw_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_psw_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_psw_s1_end_xfer <= psw_s1_end_xfer;
    end if;

  end process;

  --psw_s1_waits_for_read in a cycle, which is an e_mux
  psw_s1_waits_for_read <= psw_s1_in_a_read_cycle AND psw_s1_begins_xfer;
  --psw_s1_in_a_read_cycle assignment, which is an e_assign
  psw_s1_in_a_read_cycle <= internal_peripheral_bridge_m1_granted_psw_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= psw_s1_in_a_read_cycle;
  --psw_s1_waits_for_write in a cycle, which is an e_mux
  psw_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(psw_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --psw_s1_in_a_write_cycle assignment, which is an e_assign
  psw_s1_in_a_write_cycle <= internal_peripheral_bridge_m1_granted_psw_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= psw_s1_in_a_write_cycle;
  wait_for_psw_s1_counter <= std_logic'('0');
  --assign psw_s1_irq_from_sa = psw_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  psw_s1_irq_from_sa <= psw_s1_irq;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_granted_psw_s1 <= internal_peripheral_bridge_m1_granted_psw_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_qualified_request_psw_s1 <= internal_peripheral_bridge_m1_qualified_request_psw_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_requests_psw_s1 <= internal_peripheral_bridge_m1_requests_psw_s1;
--synthesis translate_off
    --psw/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --peripheral_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line103 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_peripheral_bridge_m1_requests_psw_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line103, now);
          write(write_line103, string'(": "));
          write(write_line103, string'("peripheral_bridge/m1 drove 0 on its 'burstcount' port while accessing slave psw/s1"));
          write(output, write_line103.all);
          deallocate (write_line103);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_nios2_fpu_burst_0_downstream_to_sdram_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_nios2_fpu_burst_0_downstream_to_sdram_s1_module;


architecture europa of rdv_fifo_for_nios2_fpu_burst_0_downstream_to_sdram_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_6;
  empty <= NOT(full_0);
  full_7 <= std_logic'('0');
  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_nios2_fpu_burst_1_downstream_to_sdram_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_nios2_fpu_burst_1_downstream_to_sdram_s1_module;


architecture europa of rdv_fifo_for_nios2_fpu_burst_1_downstream_to_sdram_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_6;
  empty <= NOT(full_0);
  full_7 <= std_logic'('0');
  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_nios2_fpu_burst_2_downstream_to_sdram_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_nios2_fpu_burst_2_downstream_to_sdram_s1_module;


architecture europa of rdv_fifo_for_nios2_fpu_burst_2_downstream_to_sdram_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_6;
  empty <= NOT(full_0);
  full_7 <= std_logic'('0');
  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_nios2_fpu_burst_3_downstream_to_sdram_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_nios2_fpu_burst_3_downstream_to_sdram_s1_module;


architecture europa of rdv_fifo_for_nios2_fpu_burst_3_downstream_to_sdram_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_6;
  empty <= NOT(full_0);
  full_7 <= std_logic'('0');
  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sdram_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_0_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal nios2_fpu_burst_0_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fpu_burst_0_downstream_latency_counter : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_1_downstream_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_1_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal nios2_fpu_burst_1_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fpu_burst_1_downstream_latency_counter : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_2_downstream_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_2_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal nios2_fpu_burst_2_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fpu_burst_2_downstream_latency_counter : IN STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_3_downstream_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal nios2_fpu_burst_3_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal nios2_fpu_burst_3_downstream_burstcount : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal nios2_fpu_burst_3_downstream_latency_counter : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_read : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_write : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_s1_readdatavalid : IN STD_LOGIC;
                 signal sdram_s1_waitrequest : IN STD_LOGIC;

              -- outputs:
                 signal d1_sdram_s1_end_xfer : OUT STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_granted_sdram_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_qualified_request_sdram_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                 signal nios2_fpu_burst_0_downstream_requests_sdram_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_granted_sdram_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_qualified_request_sdram_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                 signal nios2_fpu_burst_1_downstream_requests_sdram_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_granted_sdram_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_qualified_request_sdram_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                 signal nios2_fpu_burst_2_downstream_requests_sdram_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_granted_sdram_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_qualified_request_sdram_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                 signal nios2_fpu_burst_3_downstream_requests_sdram_s1 : OUT STD_LOGIC;
                 signal sdram_s1_address : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal sdram_s1_byteenable_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal sdram_s1_chipselect : OUT STD_LOGIC;
                 signal sdram_s1_read_n : OUT STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_s1_reset_n : OUT STD_LOGIC;
                 signal sdram_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal sdram_s1_write_n : OUT STD_LOGIC;
                 signal sdram_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity sdram_s1_arbitrator;


architecture europa of sdram_s1_arbitrator is
component rdv_fifo_for_nios2_fpu_burst_0_downstream_to_sdram_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_nios2_fpu_burst_0_downstream_to_sdram_s1_module;

component rdv_fifo_for_nios2_fpu_burst_1_downstream_to_sdram_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_nios2_fpu_burst_1_downstream_to_sdram_s1_module;

component rdv_fifo_for_nios2_fpu_burst_2_downstream_to_sdram_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_nios2_fpu_burst_2_downstream_to_sdram_s1_module;

component rdv_fifo_for_nios2_fpu_burst_3_downstream_to_sdram_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_nios2_fpu_burst_3_downstream_to_sdram_s1_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sdram_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_nios2_fpu_burst_0_downstream_granted_sdram_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_0_downstream_qualified_request_sdram_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_0_downstream_requests_sdram_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_1_downstream_granted_sdram_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_1_downstream_qualified_request_sdram_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_1_downstream_requests_sdram_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_2_downstream_granted_sdram_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_2_downstream_qualified_request_sdram_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_2_downstream_requests_sdram_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_3_downstream_granted_sdram_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_3_downstream_qualified_request_sdram_s1 :  STD_LOGIC;
                signal internal_nios2_fpu_burst_3_downstream_requests_sdram_s1 :  STD_LOGIC;
                signal internal_sdram_s1_waitrequest_from_sa :  STD_LOGIC;
                signal last_cycle_nios2_fpu_burst_0_downstream_granted_slave_sdram_s1 :  STD_LOGIC;
                signal last_cycle_nios2_fpu_burst_1_downstream_granted_slave_sdram_s1 :  STD_LOGIC;
                signal last_cycle_nios2_fpu_burst_2_downstream_granted_slave_sdram_s1 :  STD_LOGIC;
                signal last_cycle_nios2_fpu_burst_3_downstream_granted_slave_sdram_s1 :  STD_LOGIC;
                signal module_input57 :  STD_LOGIC;
                signal module_input58 :  STD_LOGIC;
                signal module_input59 :  STD_LOGIC;
                signal module_input60 :  STD_LOGIC;
                signal module_input61 :  STD_LOGIC;
                signal module_input62 :  STD_LOGIC;
                signal module_input63 :  STD_LOGIC;
                signal module_input64 :  STD_LOGIC;
                signal module_input65 :  STD_LOGIC;
                signal module_input66 :  STD_LOGIC;
                signal module_input67 :  STD_LOGIC;
                signal module_input68 :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_arbiterlock :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_arbiterlock2 :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_rdv_fifo_empty_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_rdv_fifo_output_from_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_saved_grant_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_arbiterlock :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_arbiterlock2 :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_rdv_fifo_empty_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_rdv_fifo_output_from_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_saved_grant_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_arbiterlock :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_arbiterlock2 :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_rdv_fifo_empty_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_rdv_fifo_output_from_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_saved_grant_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_arbiterlock :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_arbiterlock2 :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_continuerequest :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_rdv_fifo_empty_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_rdv_fifo_output_from_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_saved_grant_sdram_s1 :  STD_LOGIC;
                signal sdram_s1_allgrants :  STD_LOGIC;
                signal sdram_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal sdram_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sdram_s1_any_continuerequest :  STD_LOGIC;
                signal sdram_s1_arb_addend :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sdram_s1_arb_counter_enable :  STD_LOGIC;
                signal sdram_s1_arb_share_counter :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal sdram_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal sdram_s1_arb_share_set_values :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal sdram_s1_arb_winner :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sdram_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal sdram_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal sdram_s1_begins_xfer :  STD_LOGIC;
                signal sdram_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal sdram_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sdram_s1_end_xfer :  STD_LOGIC;
                signal sdram_s1_firsttransfer :  STD_LOGIC;
                signal sdram_s1_grant_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sdram_s1_in_a_read_cycle :  STD_LOGIC;
                signal sdram_s1_in_a_write_cycle :  STD_LOGIC;
                signal sdram_s1_master_qreq_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sdram_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal sdram_s1_non_bursting_master_requests :  STD_LOGIC;
                signal sdram_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal sdram_s1_reg_firsttransfer :  STD_LOGIC;
                signal sdram_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sdram_s1_slavearbiterlockenable :  STD_LOGIC;
                signal sdram_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal sdram_s1_unreg_firsttransfer :  STD_LOGIC;
                signal sdram_s1_waits_for_read :  STD_LOGIC;
                signal sdram_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_sdram_s1_from_nios2_fpu_burst_0_downstream :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal shifted_address_to_sdram_s1_from_nios2_fpu_burst_1_downstream :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal shifted_address_to_sdram_s1_from_nios2_fpu_burst_2_downstream :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal shifted_address_to_sdram_s1_from_nios2_fpu_burst_3_downstream :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_sdram_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sdram_s1_end_xfer;
    end if;

  end process;

  sdram_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((((internal_nios2_fpu_burst_0_downstream_qualified_request_sdram_s1 OR internal_nios2_fpu_burst_1_downstream_qualified_request_sdram_s1) OR internal_nios2_fpu_burst_2_downstream_qualified_request_sdram_s1) OR internal_nios2_fpu_burst_3_downstream_qualified_request_sdram_s1));
  --assign sdram_s1_readdata_from_sa = sdram_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sdram_s1_readdata_from_sa <= sdram_s1_readdata;
  internal_nios2_fpu_burst_0_downstream_requests_sdram_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_0_downstream_read OR nios2_fpu_burst_0_downstream_write)))))));
  --assign sdram_s1_waitrequest_from_sa = sdram_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_sdram_s1_waitrequest_from_sa <= sdram_s1_waitrequest;
  --assign sdram_s1_readdatavalid_from_sa = sdram_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  sdram_s1_readdatavalid_from_sa <= sdram_s1_readdatavalid;
  --sdram_s1_arb_share_counter set values, which is an e_mux
  sdram_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_0_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000") & (nios2_fpu_burst_0_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_1_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_1_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_2_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_2_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_3_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_3_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_0_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000") & (nios2_fpu_burst_0_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_1_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_1_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_2_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_2_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_3_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_3_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_0_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000") & (nios2_fpu_burst_0_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_1_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_1_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_2_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_2_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_3_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_3_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_0_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000") & (nios2_fpu_burst_0_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_1_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_1_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_2_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_2_downstream_arbitrationshare)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_3_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_3_downstream_arbitrationshare)), std_logic_vector'("00000000000000000000000000000001"))))))))))))))))), 11);
  --sdram_s1_non_bursting_master_requests mux, which is an e_mux
  sdram_s1_non_bursting_master_requests <= std_logic'('0');
  --sdram_s1_any_bursting_master_saved_grant mux, which is an e_mux
  sdram_s1_any_bursting_master_saved_grant <= ((((((((((((((nios2_fpu_burst_0_downstream_saved_grant_sdram_s1 OR nios2_fpu_burst_1_downstream_saved_grant_sdram_s1) OR nios2_fpu_burst_2_downstream_saved_grant_sdram_s1) OR nios2_fpu_burst_3_downstream_saved_grant_sdram_s1) OR nios2_fpu_burst_0_downstream_saved_grant_sdram_s1) OR nios2_fpu_burst_1_downstream_saved_grant_sdram_s1) OR nios2_fpu_burst_2_downstream_saved_grant_sdram_s1) OR nios2_fpu_burst_3_downstream_saved_grant_sdram_s1) OR nios2_fpu_burst_0_downstream_saved_grant_sdram_s1) OR nios2_fpu_burst_1_downstream_saved_grant_sdram_s1) OR nios2_fpu_burst_2_downstream_saved_grant_sdram_s1) OR nios2_fpu_burst_3_downstream_saved_grant_sdram_s1) OR nios2_fpu_burst_0_downstream_saved_grant_sdram_s1) OR nios2_fpu_burst_1_downstream_saved_grant_sdram_s1) OR nios2_fpu_burst_2_downstream_saved_grant_sdram_s1) OR nios2_fpu_burst_3_downstream_saved_grant_sdram_s1;
  --sdram_s1_arb_share_counter_next_value assignment, which is an e_assign
  sdram_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(sdram_s1_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000") & (sdram_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(sdram_s1_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000") & (sdram_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 11);
  --sdram_s1_allgrants all slave grants, which is an e_mux
  sdram_s1_allgrants <= (((((((((((((((or_reduce(sdram_s1_grant_vector)) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector));
  --sdram_s1_end_xfer assignment, which is an e_assign
  sdram_s1_end_xfer <= NOT ((sdram_s1_waits_for_read OR sdram_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_sdram_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sdram_s1 <= sdram_s1_end_xfer AND (((NOT sdram_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sdram_s1_arb_share_counter arbitration counter enable, which is an e_assign
  sdram_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sdram_s1 AND sdram_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_sdram_s1 AND NOT sdram_s1_non_bursting_master_requests));
  --sdram_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_arb_share_counter <= std_logic_vector'("00000000000");
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_s1_arb_counter_enable) = '1' then 
        sdram_s1_arb_share_counter <= sdram_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sdram_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(sdram_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_sdram_s1)) OR ((end_xfer_arb_share_counter_term_sdram_s1 AND NOT sdram_s1_non_bursting_master_requests)))) = '1' then 
        sdram_s1_slavearbiterlockenable <= or_reduce(sdram_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --nios2_fpu_burst_0/downstream sdram/s1 arbiterlock, which is an e_assign
  nios2_fpu_burst_0_downstream_arbiterlock <= sdram_s1_slavearbiterlockenable AND nios2_fpu_burst_0_downstream_continuerequest;
  --sdram_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sdram_s1_slavearbiterlockenable2 <= or_reduce(sdram_s1_arb_share_counter_next_value);
  --nios2_fpu_burst_0/downstream sdram/s1 arbiterlock2, which is an e_assign
  nios2_fpu_burst_0_downstream_arbiterlock2 <= sdram_s1_slavearbiterlockenable2 AND nios2_fpu_burst_0_downstream_continuerequest;
  --nios2_fpu_burst_1/downstream sdram/s1 arbiterlock, which is an e_assign
  nios2_fpu_burst_1_downstream_arbiterlock <= sdram_s1_slavearbiterlockenable AND nios2_fpu_burst_1_downstream_continuerequest;
  --nios2_fpu_burst_1/downstream sdram/s1 arbiterlock2, which is an e_assign
  nios2_fpu_burst_1_downstream_arbiterlock2 <= sdram_s1_slavearbiterlockenable2 AND nios2_fpu_burst_1_downstream_continuerequest;
  --nios2_fpu_burst_1/downstream granted sdram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_nios2_fpu_burst_1_downstream_granted_slave_sdram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_nios2_fpu_burst_1_downstream_granted_slave_sdram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_1_downstream_saved_grant_sdram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_s1_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_1_downstream_granted_slave_sdram_s1))))));
    end if;

  end process;

  --nios2_fpu_burst_1_downstream_continuerequest continued request, which is an e_mux
  nios2_fpu_burst_1_downstream_continuerequest <= Vector_To_Std_Logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_1_downstream_granted_slave_sdram_s1))) AND std_logic_vector'("00000000000000000000000000000001"))) OR (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_1_downstream_granted_slave_sdram_s1))) AND std_logic_vector'("00000000000000000000000000000001")))) OR (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_1_downstream_granted_slave_sdram_s1))) AND std_logic_vector'("00000000000000000000000000000001")))));
  --sdram_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  sdram_s1_any_continuerequest <= ((((((((((nios2_fpu_burst_1_downstream_continuerequest OR nios2_fpu_burst_2_downstream_continuerequest) OR nios2_fpu_burst_3_downstream_continuerequest) OR nios2_fpu_burst_0_downstream_continuerequest) OR nios2_fpu_burst_2_downstream_continuerequest) OR nios2_fpu_burst_3_downstream_continuerequest) OR nios2_fpu_burst_0_downstream_continuerequest) OR nios2_fpu_burst_1_downstream_continuerequest) OR nios2_fpu_burst_3_downstream_continuerequest) OR nios2_fpu_burst_0_downstream_continuerequest) OR nios2_fpu_burst_1_downstream_continuerequest) OR nios2_fpu_burst_2_downstream_continuerequest;
  --nios2_fpu_burst_2/downstream sdram/s1 arbiterlock, which is an e_assign
  nios2_fpu_burst_2_downstream_arbiterlock <= sdram_s1_slavearbiterlockenable AND nios2_fpu_burst_2_downstream_continuerequest;
  --nios2_fpu_burst_2/downstream sdram/s1 arbiterlock2, which is an e_assign
  nios2_fpu_burst_2_downstream_arbiterlock2 <= sdram_s1_slavearbiterlockenable2 AND nios2_fpu_burst_2_downstream_continuerequest;
  --nios2_fpu_burst_2/downstream granted sdram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_nios2_fpu_burst_2_downstream_granted_slave_sdram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_nios2_fpu_burst_2_downstream_granted_slave_sdram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_2_downstream_saved_grant_sdram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_s1_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_2_downstream_granted_slave_sdram_s1))))));
    end if;

  end process;

  --nios2_fpu_burst_2_downstream_continuerequest continued request, which is an e_mux
  nios2_fpu_burst_2_downstream_continuerequest <= Vector_To_Std_Logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_2_downstream_granted_slave_sdram_s1))) AND std_logic_vector'("00000000000000000000000000000001"))) OR (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_2_downstream_granted_slave_sdram_s1))) AND std_logic_vector'("00000000000000000000000000000001")))) OR (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_2_downstream_granted_slave_sdram_s1))) AND std_logic_vector'("00000000000000000000000000000001")))));
  --nios2_fpu_burst_3/downstream sdram/s1 arbiterlock, which is an e_assign
  nios2_fpu_burst_3_downstream_arbiterlock <= sdram_s1_slavearbiterlockenable AND nios2_fpu_burst_3_downstream_continuerequest;
  --nios2_fpu_burst_3/downstream sdram/s1 arbiterlock2, which is an e_assign
  nios2_fpu_burst_3_downstream_arbiterlock2 <= sdram_s1_slavearbiterlockenable2 AND nios2_fpu_burst_3_downstream_continuerequest;
  --nios2_fpu_burst_3/downstream granted sdram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_nios2_fpu_burst_3_downstream_granted_slave_sdram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_nios2_fpu_burst_3_downstream_granted_slave_sdram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_3_downstream_saved_grant_sdram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_s1_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_3_downstream_granted_slave_sdram_s1))))));
    end if;

  end process;

  --nios2_fpu_burst_3_downstream_continuerequest continued request, which is an e_mux
  nios2_fpu_burst_3_downstream_continuerequest <= Vector_To_Std_Logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_3_downstream_granted_slave_sdram_s1))) AND std_logic_vector'("00000000000000000000000000000001"))) OR (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_3_downstream_granted_slave_sdram_s1))) AND std_logic_vector'("00000000000000000000000000000001")))) OR (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_3_downstream_granted_slave_sdram_s1))) AND std_logic_vector'("00000000000000000000000000000001")))));
  internal_nios2_fpu_burst_0_downstream_qualified_request_sdram_s1 <= internal_nios2_fpu_burst_0_downstream_requests_sdram_s1 AND NOT ((((((nios2_fpu_burst_0_downstream_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_0_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_0_downstream_latency_counter)))))))))) OR nios2_fpu_burst_1_downstream_arbiterlock) OR nios2_fpu_burst_2_downstream_arbiterlock) OR nios2_fpu_burst_3_downstream_arbiterlock));
  --unique name for sdram_s1_move_on_to_next_transaction, which is an e_assign
  sdram_s1_move_on_to_next_transaction <= sdram_s1_readdatavalid_from_sa;
  --rdv_fifo_for_nios2_fpu_burst_0_downstream_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios2_fpu_burst_0_downstream_to_sdram_s1 : rdv_fifo_for_nios2_fpu_burst_0_downstream_to_sdram_s1_module
    port map(
      data_out => nios2_fpu_burst_0_downstream_rdv_fifo_output_from_sdram_s1,
      empty => open,
      fifo_contains_ones_n => nios2_fpu_burst_0_downstream_rdv_fifo_empty_sdram_s1,
      full => open,
      clear_fifo => module_input57,
      clk => clk,
      data_in => internal_nios2_fpu_burst_0_downstream_granted_sdram_s1,
      read => sdram_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input58,
      write => module_input59
    );

  module_input57 <= std_logic'('0');
  module_input58 <= std_logic'('0');
  module_input59 <= in_a_read_cycle AND NOT sdram_s1_waits_for_read;

  nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1_shift_register <= NOT nios2_fpu_burst_0_downstream_rdv_fifo_empty_sdram_s1;
  --local readdatavalid nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1, which is an e_mux
  nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1 <= ((sdram_s1_readdatavalid_from_sa AND nios2_fpu_burst_0_downstream_rdv_fifo_output_from_sdram_s1)) AND NOT nios2_fpu_burst_0_downstream_rdv_fifo_empty_sdram_s1;
  --sdram_s1_writedata mux, which is an e_mux
  sdram_s1_writedata <= A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_0_downstream_granted_sdram_s1)) = '1'), nios2_fpu_burst_0_downstream_writedata, A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_1_downstream_granted_sdram_s1)) = '1'), nios2_fpu_burst_1_downstream_writedata, A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_2_downstream_granted_sdram_s1)) = '1'), nios2_fpu_burst_2_downstream_writedata, nios2_fpu_burst_3_downstream_writedata)));
  internal_nios2_fpu_burst_1_downstream_requests_sdram_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_1_downstream_read OR nios2_fpu_burst_1_downstream_write)))))));
  --nios2_fpu_burst_0/downstream granted sdram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_nios2_fpu_burst_0_downstream_granted_slave_sdram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_nios2_fpu_burst_0_downstream_granted_slave_sdram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(nios2_fpu_burst_0_downstream_saved_grant_sdram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_s1_arbitration_holdoff_internal))) OR std_logic_vector'("00000000000000000000000000000000")))) /= std_logic_vector'("00000000000000000000000000000000")), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_0_downstream_granted_slave_sdram_s1))))));
    end if;

  end process;

  --nios2_fpu_burst_0_downstream_continuerequest continued request, which is an e_mux
  nios2_fpu_burst_0_downstream_continuerequest <= Vector_To_Std_Logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_0_downstream_granted_slave_sdram_s1))) AND std_logic_vector'("00000000000000000000000000000001"))) OR (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_0_downstream_granted_slave_sdram_s1))) AND std_logic_vector'("00000000000000000000000000000001")))) OR (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_nios2_fpu_burst_0_downstream_granted_slave_sdram_s1))) AND std_logic_vector'("00000000000000000000000000000001")))));
  internal_nios2_fpu_burst_1_downstream_qualified_request_sdram_s1 <= internal_nios2_fpu_burst_1_downstream_requests_sdram_s1 AND NOT ((((((nios2_fpu_burst_1_downstream_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_1_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_1_downstream_latency_counter)))))))))) OR nios2_fpu_burst_0_downstream_arbiterlock) OR nios2_fpu_burst_2_downstream_arbiterlock) OR nios2_fpu_burst_3_downstream_arbiterlock));
  --rdv_fifo_for_nios2_fpu_burst_1_downstream_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios2_fpu_burst_1_downstream_to_sdram_s1 : rdv_fifo_for_nios2_fpu_burst_1_downstream_to_sdram_s1_module
    port map(
      data_out => nios2_fpu_burst_1_downstream_rdv_fifo_output_from_sdram_s1,
      empty => open,
      fifo_contains_ones_n => nios2_fpu_burst_1_downstream_rdv_fifo_empty_sdram_s1,
      full => open,
      clear_fifo => module_input60,
      clk => clk,
      data_in => internal_nios2_fpu_burst_1_downstream_granted_sdram_s1,
      read => sdram_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input61,
      write => module_input62
    );

  module_input60 <= std_logic'('0');
  module_input61 <= std_logic'('0');
  module_input62 <= in_a_read_cycle AND NOT sdram_s1_waits_for_read;

  nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1_shift_register <= NOT nios2_fpu_burst_1_downstream_rdv_fifo_empty_sdram_s1;
  --local readdatavalid nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1, which is an e_mux
  nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1 <= ((sdram_s1_readdatavalid_from_sa AND nios2_fpu_burst_1_downstream_rdv_fifo_output_from_sdram_s1)) AND NOT nios2_fpu_burst_1_downstream_rdv_fifo_empty_sdram_s1;
  internal_nios2_fpu_burst_2_downstream_requests_sdram_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_2_downstream_read OR nios2_fpu_burst_2_downstream_write)))))));
  internal_nios2_fpu_burst_2_downstream_qualified_request_sdram_s1 <= internal_nios2_fpu_burst_2_downstream_requests_sdram_s1 AND NOT ((((((nios2_fpu_burst_2_downstream_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_2_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_2_downstream_latency_counter)))))))))) OR nios2_fpu_burst_0_downstream_arbiterlock) OR nios2_fpu_burst_1_downstream_arbiterlock) OR nios2_fpu_burst_3_downstream_arbiterlock));
  --rdv_fifo_for_nios2_fpu_burst_2_downstream_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios2_fpu_burst_2_downstream_to_sdram_s1 : rdv_fifo_for_nios2_fpu_burst_2_downstream_to_sdram_s1_module
    port map(
      data_out => nios2_fpu_burst_2_downstream_rdv_fifo_output_from_sdram_s1,
      empty => open,
      fifo_contains_ones_n => nios2_fpu_burst_2_downstream_rdv_fifo_empty_sdram_s1,
      full => open,
      clear_fifo => module_input63,
      clk => clk,
      data_in => internal_nios2_fpu_burst_2_downstream_granted_sdram_s1,
      read => sdram_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input64,
      write => module_input65
    );

  module_input63 <= std_logic'('0');
  module_input64 <= std_logic'('0');
  module_input65 <= in_a_read_cycle AND NOT sdram_s1_waits_for_read;

  nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1_shift_register <= NOT nios2_fpu_burst_2_downstream_rdv_fifo_empty_sdram_s1;
  --local readdatavalid nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1, which is an e_mux
  nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1 <= ((sdram_s1_readdatavalid_from_sa AND nios2_fpu_burst_2_downstream_rdv_fifo_output_from_sdram_s1)) AND NOT nios2_fpu_burst_2_downstream_rdv_fifo_empty_sdram_s1;
  internal_nios2_fpu_burst_3_downstream_requests_sdram_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((nios2_fpu_burst_3_downstream_read OR nios2_fpu_burst_3_downstream_write)))))));
  internal_nios2_fpu_burst_3_downstream_qualified_request_sdram_s1 <= internal_nios2_fpu_burst_3_downstream_requests_sdram_s1 AND NOT ((((((nios2_fpu_burst_3_downstream_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_3_downstream_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_3_downstream_latency_counter)))))))))) OR nios2_fpu_burst_0_downstream_arbiterlock) OR nios2_fpu_burst_1_downstream_arbiterlock) OR nios2_fpu_burst_2_downstream_arbiterlock));
  --rdv_fifo_for_nios2_fpu_burst_3_downstream_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios2_fpu_burst_3_downstream_to_sdram_s1 : rdv_fifo_for_nios2_fpu_burst_3_downstream_to_sdram_s1_module
    port map(
      data_out => nios2_fpu_burst_3_downstream_rdv_fifo_output_from_sdram_s1,
      empty => open,
      fifo_contains_ones_n => nios2_fpu_burst_3_downstream_rdv_fifo_empty_sdram_s1,
      full => open,
      clear_fifo => module_input66,
      clk => clk,
      data_in => internal_nios2_fpu_burst_3_downstream_granted_sdram_s1,
      read => sdram_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input67,
      write => module_input68
    );

  module_input66 <= std_logic'('0');
  module_input67 <= std_logic'('0');
  module_input68 <= in_a_read_cycle AND NOT sdram_s1_waits_for_read;

  nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1_shift_register <= NOT nios2_fpu_burst_3_downstream_rdv_fifo_empty_sdram_s1;
  --local readdatavalid nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1, which is an e_mux
  nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1 <= ((sdram_s1_readdatavalid_from_sa AND nios2_fpu_burst_3_downstream_rdv_fifo_output_from_sdram_s1)) AND NOT nios2_fpu_burst_3_downstream_rdv_fifo_empty_sdram_s1;
  --allow new arb cycle for sdram/s1, which is an e_assign
  sdram_s1_allow_new_arb_cycle <= ((NOT nios2_fpu_burst_0_downstream_arbiterlock AND NOT nios2_fpu_burst_1_downstream_arbiterlock) AND NOT nios2_fpu_burst_2_downstream_arbiterlock) AND NOT nios2_fpu_burst_3_downstream_arbiterlock;
  --nios2_fpu_burst_3/downstream assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  sdram_s1_master_qreq_vector(0) <= internal_nios2_fpu_burst_3_downstream_qualified_request_sdram_s1;
  --nios2_fpu_burst_3/downstream grant sdram/s1, which is an e_assign
  internal_nios2_fpu_burst_3_downstream_granted_sdram_s1 <= sdram_s1_grant_vector(0);
  --nios2_fpu_burst_3/downstream saved-grant sdram/s1, which is an e_assign
  nios2_fpu_burst_3_downstream_saved_grant_sdram_s1 <= sdram_s1_arb_winner(0);
  --nios2_fpu_burst_2/downstream assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  sdram_s1_master_qreq_vector(1) <= internal_nios2_fpu_burst_2_downstream_qualified_request_sdram_s1;
  --nios2_fpu_burst_2/downstream grant sdram/s1, which is an e_assign
  internal_nios2_fpu_burst_2_downstream_granted_sdram_s1 <= sdram_s1_grant_vector(1);
  --nios2_fpu_burst_2/downstream saved-grant sdram/s1, which is an e_assign
  nios2_fpu_burst_2_downstream_saved_grant_sdram_s1 <= sdram_s1_arb_winner(1);
  --nios2_fpu_burst_1/downstream assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  sdram_s1_master_qreq_vector(2) <= internal_nios2_fpu_burst_1_downstream_qualified_request_sdram_s1;
  --nios2_fpu_burst_1/downstream grant sdram/s1, which is an e_assign
  internal_nios2_fpu_burst_1_downstream_granted_sdram_s1 <= sdram_s1_grant_vector(2);
  --nios2_fpu_burst_1/downstream saved-grant sdram/s1, which is an e_assign
  nios2_fpu_burst_1_downstream_saved_grant_sdram_s1 <= sdram_s1_arb_winner(2);
  --nios2_fpu_burst_0/downstream assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  sdram_s1_master_qreq_vector(3) <= internal_nios2_fpu_burst_0_downstream_qualified_request_sdram_s1;
  --nios2_fpu_burst_0/downstream grant sdram/s1, which is an e_assign
  internal_nios2_fpu_burst_0_downstream_granted_sdram_s1 <= sdram_s1_grant_vector(3);
  --nios2_fpu_burst_0/downstream saved-grant sdram/s1, which is an e_assign
  nios2_fpu_burst_0_downstream_saved_grant_sdram_s1 <= sdram_s1_arb_winner(3);
  --sdram/s1 chosen-master double-vector, which is an e_assign
  sdram_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((sdram_s1_master_qreq_vector & sdram_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT sdram_s1_master_qreq_vector & NOT sdram_s1_master_qreq_vector))) + (std_logic_vector'("00000") & (sdram_s1_arb_addend))))), 8);
  --stable onehot encoding of arb winner
  sdram_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((sdram_s1_allow_new_arb_cycle AND or_reduce(sdram_s1_grant_vector)))) = '1'), sdram_s1_grant_vector, sdram_s1_saved_chosen_master_vector);
  --saved sdram_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_saved_chosen_master_vector <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_s1_allow_new_arb_cycle) = '1' then 
        sdram_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(sdram_s1_grant_vector)) = '1'), sdram_s1_grant_vector, sdram_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  sdram_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((sdram_s1_chosen_master_double_vector(3) OR sdram_s1_chosen_master_double_vector(7)))) & A_ToStdLogicVector(((sdram_s1_chosen_master_double_vector(2) OR sdram_s1_chosen_master_double_vector(6)))) & A_ToStdLogicVector(((sdram_s1_chosen_master_double_vector(1) OR sdram_s1_chosen_master_double_vector(5)))) & A_ToStdLogicVector(((sdram_s1_chosen_master_double_vector(0) OR sdram_s1_chosen_master_double_vector(4)))));
  --sdram/s1 chosen master rotated left, which is an e_assign
  sdram_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(sdram_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("0000")), (std_logic_vector'("0000000000000000000000000000") & ((A_SLL(sdram_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 4);
  --sdram/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_arb_addend <= std_logic_vector'("0001");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(sdram_s1_grant_vector)) = '1' then 
        sdram_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(sdram_s1_end_xfer) = '1'), sdram_s1_chosen_master_rot_left, sdram_s1_grant_vector);
      end if;
    end if;

  end process;

  --sdram_s1_reset_n assignment, which is an e_assign
  sdram_s1_reset_n <= reset_n;
  sdram_s1_chipselect <= ((internal_nios2_fpu_burst_0_downstream_granted_sdram_s1 OR internal_nios2_fpu_burst_1_downstream_granted_sdram_s1) OR internal_nios2_fpu_burst_2_downstream_granted_sdram_s1) OR internal_nios2_fpu_burst_3_downstream_granted_sdram_s1;
  --sdram_s1_firsttransfer first transaction, which is an e_assign
  sdram_s1_firsttransfer <= A_WE_StdLogic((std_logic'(sdram_s1_begins_xfer) = '1'), sdram_s1_unreg_firsttransfer, sdram_s1_reg_firsttransfer);
  --sdram_s1_unreg_firsttransfer first transaction, which is an e_assign
  sdram_s1_unreg_firsttransfer <= NOT ((sdram_s1_slavearbiterlockenable AND sdram_s1_any_continuerequest));
  --sdram_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_s1_begins_xfer) = '1' then 
        sdram_s1_reg_firsttransfer <= sdram_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sdram_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sdram_s1_beginbursttransfer_internal <= sdram_s1_begins_xfer;
  --sdram_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  sdram_s1_arbitration_holdoff_internal <= sdram_s1_begins_xfer AND sdram_s1_firsttransfer;
  --~sdram_s1_read_n assignment, which is an e_mux
  sdram_s1_read_n <= NOT ((((((internal_nios2_fpu_burst_0_downstream_granted_sdram_s1 AND nios2_fpu_burst_0_downstream_read)) OR ((internal_nios2_fpu_burst_1_downstream_granted_sdram_s1 AND nios2_fpu_burst_1_downstream_read))) OR ((internal_nios2_fpu_burst_2_downstream_granted_sdram_s1 AND nios2_fpu_burst_2_downstream_read))) OR ((internal_nios2_fpu_burst_3_downstream_granted_sdram_s1 AND nios2_fpu_burst_3_downstream_read))));
  --~sdram_s1_write_n assignment, which is an e_mux
  sdram_s1_write_n <= NOT ((((((internal_nios2_fpu_burst_0_downstream_granted_sdram_s1 AND nios2_fpu_burst_0_downstream_write)) OR ((internal_nios2_fpu_burst_1_downstream_granted_sdram_s1 AND nios2_fpu_burst_1_downstream_write))) OR ((internal_nios2_fpu_burst_2_downstream_granted_sdram_s1 AND nios2_fpu_burst_2_downstream_write))) OR ((internal_nios2_fpu_burst_3_downstream_granted_sdram_s1 AND nios2_fpu_burst_3_downstream_write))));
  shifted_address_to_sdram_s1_from_nios2_fpu_burst_0_downstream <= nios2_fpu_burst_0_downstream_address_to_slave;
  --sdram_s1_address mux, which is an e_mux
  sdram_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_0_downstream_granted_sdram_s1)) = '1'), (A_SRL(shifted_address_to_sdram_s1_from_nios2_fpu_burst_0_downstream,std_logic_vector'("00000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_1_downstream_granted_sdram_s1)) = '1'), (A_SRL(shifted_address_to_sdram_s1_from_nios2_fpu_burst_1_downstream,std_logic_vector'("00000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_2_downstream_granted_sdram_s1)) = '1'), (A_SRL(shifted_address_to_sdram_s1_from_nios2_fpu_burst_2_downstream,std_logic_vector'("00000000000000000000000000000001"))), (A_SRL(shifted_address_to_sdram_s1_from_nios2_fpu_burst_3_downstream,std_logic_vector'("00000000000000000000000000000001")))))), 24);
  shifted_address_to_sdram_s1_from_nios2_fpu_burst_1_downstream <= nios2_fpu_burst_1_downstream_address_to_slave;
  shifted_address_to_sdram_s1_from_nios2_fpu_burst_2_downstream <= nios2_fpu_burst_2_downstream_address_to_slave;
  shifted_address_to_sdram_s1_from_nios2_fpu_burst_3_downstream <= nios2_fpu_burst_3_downstream_address_to_slave;
  --d1_sdram_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sdram_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sdram_s1_end_xfer <= sdram_s1_end_xfer;
    end if;

  end process;

  --sdram_s1_waits_for_read in a cycle, which is an e_mux
  sdram_s1_waits_for_read <= sdram_s1_in_a_read_cycle AND internal_sdram_s1_waitrequest_from_sa;
  --sdram_s1_in_a_read_cycle assignment, which is an e_assign
  sdram_s1_in_a_read_cycle <= ((((internal_nios2_fpu_burst_0_downstream_granted_sdram_s1 AND nios2_fpu_burst_0_downstream_read)) OR ((internal_nios2_fpu_burst_1_downstream_granted_sdram_s1 AND nios2_fpu_burst_1_downstream_read))) OR ((internal_nios2_fpu_burst_2_downstream_granted_sdram_s1 AND nios2_fpu_burst_2_downstream_read))) OR ((internal_nios2_fpu_burst_3_downstream_granted_sdram_s1 AND nios2_fpu_burst_3_downstream_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sdram_s1_in_a_read_cycle;
  --sdram_s1_waits_for_write in a cycle, which is an e_mux
  sdram_s1_waits_for_write <= sdram_s1_in_a_write_cycle AND internal_sdram_s1_waitrequest_from_sa;
  --sdram_s1_in_a_write_cycle assignment, which is an e_assign
  sdram_s1_in_a_write_cycle <= ((((internal_nios2_fpu_burst_0_downstream_granted_sdram_s1 AND nios2_fpu_burst_0_downstream_write)) OR ((internal_nios2_fpu_burst_1_downstream_granted_sdram_s1 AND nios2_fpu_burst_1_downstream_write))) OR ((internal_nios2_fpu_burst_2_downstream_granted_sdram_s1 AND nios2_fpu_burst_2_downstream_write))) OR ((internal_nios2_fpu_burst_3_downstream_granted_sdram_s1 AND nios2_fpu_burst_3_downstream_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sdram_s1_in_a_write_cycle;
  wait_for_sdram_s1_counter <= std_logic'('0');
  --~sdram_s1_byteenable_n byte enable port mux, which is an e_mux
  sdram_s1_byteenable_n <= A_EXT (NOT (A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_0_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (nios2_fpu_burst_0_downstream_byteenable)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_1_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (nios2_fpu_burst_1_downstream_byteenable)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_2_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (nios2_fpu_burst_2_downstream_byteenable)), A_WE_StdLogicVector((std_logic'((internal_nios2_fpu_burst_3_downstream_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (nios2_fpu_burst_3_downstream_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))))))), 2);
  --vhdl renameroo for output signals
  nios2_fpu_burst_0_downstream_granted_sdram_s1 <= internal_nios2_fpu_burst_0_downstream_granted_sdram_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_0_downstream_qualified_request_sdram_s1 <= internal_nios2_fpu_burst_0_downstream_qualified_request_sdram_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_0_downstream_requests_sdram_s1 <= internal_nios2_fpu_burst_0_downstream_requests_sdram_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_1_downstream_granted_sdram_s1 <= internal_nios2_fpu_burst_1_downstream_granted_sdram_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_1_downstream_qualified_request_sdram_s1 <= internal_nios2_fpu_burst_1_downstream_qualified_request_sdram_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_1_downstream_requests_sdram_s1 <= internal_nios2_fpu_burst_1_downstream_requests_sdram_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_2_downstream_granted_sdram_s1 <= internal_nios2_fpu_burst_2_downstream_granted_sdram_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_2_downstream_qualified_request_sdram_s1 <= internal_nios2_fpu_burst_2_downstream_qualified_request_sdram_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_2_downstream_requests_sdram_s1 <= internal_nios2_fpu_burst_2_downstream_requests_sdram_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_3_downstream_granted_sdram_s1 <= internal_nios2_fpu_burst_3_downstream_granted_sdram_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_3_downstream_qualified_request_sdram_s1 <= internal_nios2_fpu_burst_3_downstream_qualified_request_sdram_s1;
  --vhdl renameroo for output signals
  nios2_fpu_burst_3_downstream_requests_sdram_s1 <= internal_nios2_fpu_burst_3_downstream_requests_sdram_s1;
  --vhdl renameroo for output signals
  sdram_s1_waitrequest_from_sa <= internal_sdram_s1_waitrequest_from_sa;
--synthesis translate_off
    --sdram/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --nios2_fpu_burst_0/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line104 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_0_downstream_requests_sdram_s1 AND to_std_logic((((std_logic_vector'("000000000000000000000") & (nios2_fpu_burst_0_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line104, now);
          write(write_line104, string'(": "));
          write(write_line104, string'("nios2_fpu_burst_0/downstream drove 0 on its 'arbitrationshare' port while accessing slave sdram/s1"));
          write(output, write_line104.all);
          deallocate (write_line104);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_0/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line105 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_0_downstream_requests_sdram_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_0_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line105, now);
          write(write_line105, string'(": "));
          write(write_line105, string'("nios2_fpu_burst_0/downstream drove 0 on its 'burstcount' port while accessing slave sdram/s1"));
          write(output, write_line105.all);
          deallocate (write_line105);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_1/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line106 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_1_downstream_requests_sdram_s1 AND to_std_logic((((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_1_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line106, now);
          write(write_line106, string'(": "));
          write(write_line106, string'("nios2_fpu_burst_1/downstream drove 0 on its 'arbitrationshare' port while accessing slave sdram/s1"));
          write(output, write_line106.all);
          deallocate (write_line106);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_1/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line107 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_1_downstream_requests_sdram_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_1_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line107, now);
          write(write_line107, string'(": "));
          write(write_line107, string'("nios2_fpu_burst_1/downstream drove 0 on its 'burstcount' port while accessing slave sdram/s1"));
          write(output, write_line107.all);
          deallocate (write_line107);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_2/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line108 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_2_downstream_requests_sdram_s1 AND to_std_logic((((std_logic_vector'("000000000000000000000000000") & (nios2_fpu_burst_2_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line108, now);
          write(write_line108, string'(": "));
          write(write_line108, string'("nios2_fpu_burst_2/downstream drove 0 on its 'arbitrationshare' port while accessing slave sdram/s1"));
          write(output, write_line108.all);
          deallocate (write_line108);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_2/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line109 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_2_downstream_requests_sdram_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_2_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line109, now);
          write(write_line109, string'(": "));
          write(write_line109, string'("nios2_fpu_burst_2/downstream drove 0 on its 'burstcount' port while accessing slave sdram/s1"));
          write(output, write_line109.all);
          deallocate (write_line109);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_3/downstream non-zero arbitrationshare assertion, which is an e_process
    process (clk)
    VARIABLE write_line110 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_3_downstream_requests_sdram_s1 AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (nios2_fpu_burst_3_downstream_arbitrationshare)) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line110, now);
          write(write_line110, string'(": "));
          write(write_line110, string'("nios2_fpu_burst_3/downstream drove 0 on its 'arbitrationshare' port while accessing slave sdram/s1"));
          write(output, write_line110.all);
          deallocate (write_line110);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --nios2_fpu_burst_3/downstream non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line111 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_nios2_fpu_burst_3_downstream_requests_sdram_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_3_downstream_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line111, now);
          write(write_line111, string'(": "));
          write(write_line111, string'("nios2_fpu_burst_3/downstream drove 0 on its 'burstcount' port while accessing slave sdram/s1"));
          write(output, write_line111.all);
          deallocate (write_line111);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line112 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("0000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_0_downstream_granted_sdram_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_1_downstream_granted_sdram_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_2_downstream_granted_sdram_s1)))))) + (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(internal_nios2_fpu_burst_3_downstream_granted_sdram_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line112, now);
          write(write_line112, string'(": "));
          write(write_line112, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line112.all);
          deallocate (write_line112);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line113 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("0000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_0_downstream_saved_grant_sdram_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_1_downstream_saved_grant_sdram_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_2_downstream_saved_grant_sdram_s1)))))) + (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(nios2_fpu_burst_3_downstream_saved_grant_sdram_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line113, now);
          write(write_line113, string'(": "));
          write(write_line113, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line113.all);
          deallocate (write_line113);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity spu_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                 signal peripheral_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                 signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read : IN STD_LOGIC;
                 signal peripheral_bridge_m1_write : IN STD_LOGIC;
                 signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal spu_s1_irq : IN STD_LOGIC;
                 signal spu_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal spu_s1_waitrequest : IN STD_LOGIC;

              -- outputs:
                 signal d1_spu_s1_end_xfer : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_granted_spu_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_spu_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_spu_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_requests_spu_s1 : OUT STD_LOGIC;
                 signal spu_s1_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                 signal spu_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal spu_s1_chipselect : OUT STD_LOGIC;
                 signal spu_s1_irq_from_sa : OUT STD_LOGIC;
                 signal spu_s1_read : OUT STD_LOGIC;
                 signal spu_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal spu_s1_reset : OUT STD_LOGIC;
                 signal spu_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal spu_s1_write : OUT STD_LOGIC;
                 signal spu_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity spu_s1_arbitrator;


architecture europa of spu_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_spu_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_granted_spu_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_qualified_request_spu_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_requests_spu_s1 :  STD_LOGIC;
                signal internal_spu_s1_waitrequest_from_sa :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal peripheral_bridge_m1_continuerequest :  STD_LOGIC;
                signal peripheral_bridge_m1_saved_grant_spu_s1 :  STD_LOGIC;
                signal shifted_address_to_spu_s1_from_peripheral_bridge_m1 :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal spu_s1_allgrants :  STD_LOGIC;
                signal spu_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal spu_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal spu_s1_any_continuerequest :  STD_LOGIC;
                signal spu_s1_arb_counter_enable :  STD_LOGIC;
                signal spu_s1_arb_share_counter :  STD_LOGIC;
                signal spu_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal spu_s1_arb_share_set_values :  STD_LOGIC;
                signal spu_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal spu_s1_begins_xfer :  STD_LOGIC;
                signal spu_s1_end_xfer :  STD_LOGIC;
                signal spu_s1_firsttransfer :  STD_LOGIC;
                signal spu_s1_grant_vector :  STD_LOGIC;
                signal spu_s1_in_a_read_cycle :  STD_LOGIC;
                signal spu_s1_in_a_write_cycle :  STD_LOGIC;
                signal spu_s1_master_qreq_vector :  STD_LOGIC;
                signal spu_s1_non_bursting_master_requests :  STD_LOGIC;
                signal spu_s1_reg_firsttransfer :  STD_LOGIC;
                signal spu_s1_slavearbiterlockenable :  STD_LOGIC;
                signal spu_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal spu_s1_unreg_firsttransfer :  STD_LOGIC;
                signal spu_s1_waits_for_read :  STD_LOGIC;
                signal spu_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_spu_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT spu_s1_end_xfer;
    end if;

  end process;

  spu_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_peripheral_bridge_m1_qualified_request_spu_s1);
  --assign spu_s1_readdata_from_sa = spu_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  spu_s1_readdata_from_sa <= spu_s1_readdata;
  internal_peripheral_bridge_m1_requests_spu_s1 <= to_std_logic(((Std_Logic_Vector'(peripheral_bridge_m1_address_to_slave(12 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("1000000000000")))) AND peripheral_bridge_m1_chipselect;
  --assign spu_s1_waitrequest_from_sa = spu_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_spu_s1_waitrequest_from_sa <= spu_s1_waitrequest;
  --spu_s1_arb_share_counter set values, which is an e_mux
  spu_s1_arb_share_set_values <= std_logic'('1');
  --spu_s1_non_bursting_master_requests mux, which is an e_mux
  spu_s1_non_bursting_master_requests <= internal_peripheral_bridge_m1_requests_spu_s1;
  --spu_s1_any_bursting_master_saved_grant mux, which is an e_mux
  spu_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --spu_s1_arb_share_counter_next_value assignment, which is an e_assign
  spu_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(spu_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(spu_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(spu_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(spu_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --spu_s1_allgrants all slave grants, which is an e_mux
  spu_s1_allgrants <= spu_s1_grant_vector;
  --spu_s1_end_xfer assignment, which is an e_assign
  spu_s1_end_xfer <= NOT ((spu_s1_waits_for_read OR spu_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_spu_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_spu_s1 <= spu_s1_end_xfer AND (((NOT spu_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --spu_s1_arb_share_counter arbitration counter enable, which is an e_assign
  spu_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_spu_s1 AND spu_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_spu_s1 AND NOT spu_s1_non_bursting_master_requests));
  --spu_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      spu_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(spu_s1_arb_counter_enable) = '1' then 
        spu_s1_arb_share_counter <= spu_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --spu_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      spu_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((spu_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_spu_s1)) OR ((end_xfer_arb_share_counter_term_spu_s1 AND NOT spu_s1_non_bursting_master_requests)))) = '1' then 
        spu_s1_slavearbiterlockenable <= spu_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --peripheral_bridge/m1 spu/s1 arbiterlock, which is an e_assign
  peripheral_bridge_m1_arbiterlock <= spu_s1_slavearbiterlockenable AND peripheral_bridge_m1_continuerequest;
  --spu_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  spu_s1_slavearbiterlockenable2 <= spu_s1_arb_share_counter_next_value;
  --peripheral_bridge/m1 spu/s1 arbiterlock2, which is an e_assign
  peripheral_bridge_m1_arbiterlock2 <= spu_s1_slavearbiterlockenable2 AND peripheral_bridge_m1_continuerequest;
  --spu_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  spu_s1_any_continuerequest <= std_logic'('1');
  --peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  peripheral_bridge_m1_continuerequest <= std_logic'('1');
  internal_peripheral_bridge_m1_qualified_request_spu_s1 <= internal_peripheral_bridge_m1_requests_spu_s1 AND NOT ((((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid peripheral_bridge_m1_read_data_valid_spu_s1, which is an e_mux
  peripheral_bridge_m1_read_data_valid_spu_s1 <= (internal_peripheral_bridge_m1_granted_spu_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect))) AND NOT spu_s1_waits_for_read;
  --spu_s1_writedata mux, which is an e_mux
  spu_s1_writedata <= peripheral_bridge_m1_writedata;
  --master is always granted when requested
  internal_peripheral_bridge_m1_granted_spu_s1 <= internal_peripheral_bridge_m1_qualified_request_spu_s1;
  --peripheral_bridge/m1 saved-grant spu/s1, which is an e_assign
  peripheral_bridge_m1_saved_grant_spu_s1 <= internal_peripheral_bridge_m1_requests_spu_s1;
  --allow new arb cycle for spu/s1, which is an e_assign
  spu_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  spu_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  spu_s1_master_qreq_vector <= std_logic'('1');
  --~spu_s1_reset assignment, which is an e_assign
  spu_s1_reset <= NOT reset_n;
  spu_s1_chipselect <= internal_peripheral_bridge_m1_granted_spu_s1;
  --spu_s1_firsttransfer first transaction, which is an e_assign
  spu_s1_firsttransfer <= A_WE_StdLogic((std_logic'(spu_s1_begins_xfer) = '1'), spu_s1_unreg_firsttransfer, spu_s1_reg_firsttransfer);
  --spu_s1_unreg_firsttransfer first transaction, which is an e_assign
  spu_s1_unreg_firsttransfer <= NOT ((spu_s1_slavearbiterlockenable AND spu_s1_any_continuerequest));
  --spu_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      spu_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(spu_s1_begins_xfer) = '1' then 
        spu_s1_reg_firsttransfer <= spu_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --spu_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  spu_s1_beginbursttransfer_internal <= spu_s1_begins_xfer;
  --spu_s1_read assignment, which is an e_mux
  spu_s1_read <= internal_peripheral_bridge_m1_granted_spu_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --spu_s1_write assignment, which is an e_mux
  spu_s1_write <= internal_peripheral_bridge_m1_granted_spu_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect));
  shifted_address_to_spu_s1_from_peripheral_bridge_m1 <= peripheral_bridge_m1_address_to_slave;
  --spu_s1_address mux, which is an e_mux
  spu_s1_address <= A_EXT (A_SRL(shifted_address_to_spu_s1_from_peripheral_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 9);
  --d1_spu_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_spu_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_spu_s1_end_xfer <= spu_s1_end_xfer;
    end if;

  end process;

  --spu_s1_waits_for_read in a cycle, which is an e_mux
  spu_s1_waits_for_read <= spu_s1_in_a_read_cycle AND internal_spu_s1_waitrequest_from_sa;
  --spu_s1_in_a_read_cycle assignment, which is an e_assign
  spu_s1_in_a_read_cycle <= internal_peripheral_bridge_m1_granted_spu_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= spu_s1_in_a_read_cycle;
  --spu_s1_waits_for_write in a cycle, which is an e_mux
  spu_s1_waits_for_write <= spu_s1_in_a_write_cycle AND internal_spu_s1_waitrequest_from_sa;
  --spu_s1_in_a_write_cycle assignment, which is an e_assign
  spu_s1_in_a_write_cycle <= internal_peripheral_bridge_m1_granted_spu_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= spu_s1_in_a_write_cycle;
  wait_for_spu_s1_counter <= std_logic'('0');
  --spu_s1_byteenable byte enable port mux, which is an e_mux
  spu_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_peripheral_bridge_m1_granted_spu_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (peripheral_bridge_m1_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --assign spu_s1_irq_from_sa = spu_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  spu_s1_irq_from_sa <= spu_s1_irq;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_granted_spu_s1 <= internal_peripheral_bridge_m1_granted_spu_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_qualified_request_spu_s1 <= internal_peripheral_bridge_m1_qualified_request_spu_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_requests_spu_s1 <= internal_peripheral_bridge_m1_requests_spu_s1;
  --vhdl renameroo for output signals
  spu_s1_waitrequest_from_sa <= internal_spu_s1_waitrequest_from_sa;
--synthesis translate_off
    --spu/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --peripheral_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line114 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_peripheral_bridge_m1_requests_spu_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line114, now);
          write(write_line114, string'(": "));
          write(write_line114, string'("peripheral_bridge/m1 drove 0 on its 'burstcount' port while accessing slave spu/s1"));
          write(output, write_line114.all);
          deallocate (write_line114);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity spu_m1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_nios2_fpu_burst_3_upstream_end_xfer : IN STD_LOGIC;
                 signal nios2_fpu_burst_3_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_3_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal spu_m1_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal spu_m1_burstcount : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal spu_m1_granted_nios2_fpu_burst_3_upstream : IN STD_LOGIC;
                 signal spu_m1_qualified_request_nios2_fpu_burst_3_upstream : IN STD_LOGIC;
                 signal spu_m1_read : IN STD_LOGIC;
                 signal spu_m1_read_data_valid_nios2_fpu_burst_3_upstream : IN STD_LOGIC;
                 signal spu_m1_read_data_valid_nios2_fpu_burst_3_upstream_shift_register : IN STD_LOGIC;
                 signal spu_m1_requests_nios2_fpu_burst_3_upstream : IN STD_LOGIC;

              -- outputs:
                 signal spu_m1_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal spu_m1_latency_counter : OUT STD_LOGIC;
                 signal spu_m1_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal spu_m1_readdatavalid : OUT STD_LOGIC;
                 signal spu_m1_waitrequest : OUT STD_LOGIC
              );
end entity spu_m1_arbitrator;


architecture europa of spu_m1_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_spu_m1_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal internal_spu_m1_waitrequest :  STD_LOGIC;
                signal pre_flush_spu_m1_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal spu_m1_address_last_time :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal spu_m1_burstcount_last_time :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal spu_m1_read_last_time :  STD_LOGIC;
                signal spu_m1_run :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((spu_m1_qualified_request_nios2_fpu_burst_3_upstream OR NOT spu_m1_requests_nios2_fpu_burst_3_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT spu_m1_qualified_request_nios2_fpu_burst_3_upstream OR NOT (spu_m1_read))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_3_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((spu_m1_read))))))))));
  --cascaded wait assignment, which is an e_assign
  spu_m1_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_spu_m1_address_to_slave <= spu_m1_address(24 DOWNTO 0);
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_spu_m1_readdatavalid <= spu_m1_read_data_valid_nios2_fpu_burst_3_upstream;
  --latent slave read data valid which is not flushed, which is an e_mux
  spu_m1_readdatavalid <= Vector_To_Std_Logic((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_spu_m1_readdatavalid)))));
  --spu/m1 readdata mux, which is an e_mux
  spu_m1_readdata <= nios2_fpu_burst_3_upstream_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_spu_m1_waitrequest <= NOT spu_m1_run;
  --latent max counter, which is an e_assign
  spu_m1_latency_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  spu_m1_address_to_slave <= internal_spu_m1_address_to_slave;
  --vhdl renameroo for output signals
  spu_m1_waitrequest <= internal_spu_m1_waitrequest;
--synthesis translate_off
    --spu_m1_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        spu_m1_address_last_time <= std_logic_vector'("0000000000000000000000000");
      elsif clk'event and clk = '1' then
        spu_m1_address_last_time <= spu_m1_address;
      end if;

    end process;

    --spu/m1 waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_spu_m1_waitrequest AND (spu_m1_read);
      end if;

    end process;

    --spu_m1_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line115 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((spu_m1_address /= spu_m1_address_last_time))))) = '1' then 
          write(write_line115, now);
          write(write_line115, string'(": "));
          write(write_line115, string'("spu_m1_address did not heed wait!!!"));
          write(output, write_line115.all);
          deallocate (write_line115);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --spu_m1_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        spu_m1_burstcount_last_time <= std_logic_vector'("000");
      elsif clk'event and clk = '1' then
        spu_m1_burstcount_last_time <= spu_m1_burstcount;
      end if;

    end process;

    --spu_m1_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line116 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((spu_m1_burstcount /= spu_m1_burstcount_last_time))))) = '1' then 
          write(write_line116, now);
          write(write_line116, string'(": "));
          write(write_line116, string'("spu_m1_burstcount did not heed wait!!!"));
          write(output, write_line116.all);
          deallocate (write_line116);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --spu_m1_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        spu_m1_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        spu_m1_read_last_time <= spu_m1_read;
      end if;

    end process;

    --spu_m1_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line117 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(spu_m1_read) /= std_logic'(spu_m1_read_last_time)))))) = '1' then 
          write(write_line117, now);
          write(write_line117, string'(": "));
          write(write_line117, string'("spu_m1_read did not heed wait!!!"));
          write(output, write_line117.all);
          deallocate (write_line117);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sysid_control_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                 signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                 signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read : IN STD_LOGIC;
                 signal peripheral_bridge_m1_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sysid_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal d1_sysid_control_slave_end_xfer : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_granted_sysid_control_slave : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_sysid_control_slave : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_sysid_control_slave : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_requests_sysid_control_slave : OUT STD_LOGIC;
                 signal sysid_control_slave_address : OUT STD_LOGIC;
                 signal sysid_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sysid_control_slave_reset_n : OUT STD_LOGIC
              );
end entity sysid_control_slave_arbitrator;


architecture europa of sysid_control_slave_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sysid_control_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_granted_sysid_control_slave :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_qualified_request_sysid_control_slave :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_requests_sysid_control_slave :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal peripheral_bridge_m1_continuerequest :  STD_LOGIC;
                signal peripheral_bridge_m1_saved_grant_sysid_control_slave :  STD_LOGIC;
                signal shifted_address_to_sysid_control_slave_from_peripheral_bridge_m1 :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal sysid_control_slave_allgrants :  STD_LOGIC;
                signal sysid_control_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal sysid_control_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sysid_control_slave_any_continuerequest :  STD_LOGIC;
                signal sysid_control_slave_arb_counter_enable :  STD_LOGIC;
                signal sysid_control_slave_arb_share_counter :  STD_LOGIC;
                signal sysid_control_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal sysid_control_slave_arb_share_set_values :  STD_LOGIC;
                signal sysid_control_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal sysid_control_slave_begins_xfer :  STD_LOGIC;
                signal sysid_control_slave_end_xfer :  STD_LOGIC;
                signal sysid_control_slave_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_grant_vector :  STD_LOGIC;
                signal sysid_control_slave_in_a_read_cycle :  STD_LOGIC;
                signal sysid_control_slave_in_a_write_cycle :  STD_LOGIC;
                signal sysid_control_slave_master_qreq_vector :  STD_LOGIC;
                signal sysid_control_slave_non_bursting_master_requests :  STD_LOGIC;
                signal sysid_control_slave_reg_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_slavearbiterlockenable :  STD_LOGIC;
                signal sysid_control_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal sysid_control_slave_unreg_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_waits_for_read :  STD_LOGIC;
                signal sysid_control_slave_waits_for_write :  STD_LOGIC;
                signal wait_for_sysid_control_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sysid_control_slave_end_xfer;
    end if;

  end process;

  sysid_control_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_peripheral_bridge_m1_qualified_request_sysid_control_slave);
  --assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sysid_control_slave_readdata_from_sa <= sysid_control_slave_readdata;
  internal_peripheral_bridge_m1_requests_sysid_control_slave <= ((to_std_logic(((Std_Logic_Vector'(peripheral_bridge_m1_address_to_slave(12 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("0000000000000")))) AND peripheral_bridge_m1_chipselect)) AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --sysid_control_slave_arb_share_counter set values, which is an e_mux
  sysid_control_slave_arb_share_set_values <= std_logic'('1');
  --sysid_control_slave_non_bursting_master_requests mux, which is an e_mux
  sysid_control_slave_non_bursting_master_requests <= internal_peripheral_bridge_m1_requests_sysid_control_slave;
  --sysid_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  sysid_control_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --sysid_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  sysid_control_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sysid_control_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysid_control_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(sysid_control_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysid_control_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --sysid_control_slave_allgrants all slave grants, which is an e_mux
  sysid_control_slave_allgrants <= sysid_control_slave_grant_vector;
  --sysid_control_slave_end_xfer assignment, which is an e_assign
  sysid_control_slave_end_xfer <= NOT ((sysid_control_slave_waits_for_read OR sysid_control_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_sysid_control_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sysid_control_slave <= sysid_control_slave_end_xfer AND (((NOT sysid_control_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sysid_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  sysid_control_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sysid_control_slave AND sysid_control_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_sysid_control_slave AND NOT sysid_control_slave_non_bursting_master_requests));
  --sysid_control_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(sysid_control_slave_arb_counter_enable) = '1' then 
        sysid_control_slave_arb_share_counter <= sysid_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sysid_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sysid_control_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_sysid_control_slave)) OR ((end_xfer_arb_share_counter_term_sysid_control_slave AND NOT sysid_control_slave_non_bursting_master_requests)))) = '1' then 
        sysid_control_slave_slavearbiterlockenable <= sysid_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --peripheral_bridge/m1 sysid/control_slave arbiterlock, which is an e_assign
  peripheral_bridge_m1_arbiterlock <= sysid_control_slave_slavearbiterlockenable AND peripheral_bridge_m1_continuerequest;
  --sysid_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sysid_control_slave_slavearbiterlockenable2 <= sysid_control_slave_arb_share_counter_next_value;
  --peripheral_bridge/m1 sysid/control_slave arbiterlock2, which is an e_assign
  peripheral_bridge_m1_arbiterlock2 <= sysid_control_slave_slavearbiterlockenable2 AND peripheral_bridge_m1_continuerequest;
  --sysid_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  sysid_control_slave_any_continuerequest <= std_logic'('1');
  --peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  peripheral_bridge_m1_continuerequest <= std_logic'('1');
  internal_peripheral_bridge_m1_qualified_request_sysid_control_slave <= internal_peripheral_bridge_m1_requests_sysid_control_slave AND NOT ((((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid peripheral_bridge_m1_read_data_valid_sysid_control_slave, which is an e_mux
  peripheral_bridge_m1_read_data_valid_sysid_control_slave <= (internal_peripheral_bridge_m1_granted_sysid_control_slave AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect))) AND NOT sysid_control_slave_waits_for_read;
  --master is always granted when requested
  internal_peripheral_bridge_m1_granted_sysid_control_slave <= internal_peripheral_bridge_m1_qualified_request_sysid_control_slave;
  --peripheral_bridge/m1 saved-grant sysid/control_slave, which is an e_assign
  peripheral_bridge_m1_saved_grant_sysid_control_slave <= internal_peripheral_bridge_m1_requests_sysid_control_slave;
  --allow new arb cycle for sysid/control_slave, which is an e_assign
  sysid_control_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sysid_control_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sysid_control_slave_master_qreq_vector <= std_logic'('1');
  --sysid_control_slave_reset_n assignment, which is an e_assign
  sysid_control_slave_reset_n <= reset_n;
  --sysid_control_slave_firsttransfer first transaction, which is an e_assign
  sysid_control_slave_firsttransfer <= A_WE_StdLogic((std_logic'(sysid_control_slave_begins_xfer) = '1'), sysid_control_slave_unreg_firsttransfer, sysid_control_slave_reg_firsttransfer);
  --sysid_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  sysid_control_slave_unreg_firsttransfer <= NOT ((sysid_control_slave_slavearbiterlockenable AND sysid_control_slave_any_continuerequest));
  --sysid_control_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sysid_control_slave_begins_xfer) = '1' then 
        sysid_control_slave_reg_firsttransfer <= sysid_control_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sysid_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sysid_control_slave_beginbursttransfer_internal <= sysid_control_slave_begins_xfer;
  shifted_address_to_sysid_control_slave_from_peripheral_bridge_m1 <= peripheral_bridge_m1_address_to_slave;
  --sysid_control_slave_address mux, which is an e_mux
  sysid_control_slave_address <= Vector_To_Std_Logic(A_SRL(shifted_address_to_sysid_control_slave_from_peripheral_bridge_m1,std_logic_vector'("00000000000000000000000000000010")));
  --d1_sysid_control_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sysid_control_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sysid_control_slave_end_xfer <= sysid_control_slave_end_xfer;
    end if;

  end process;

  --sysid_control_slave_waits_for_read in a cycle, which is an e_mux
  sysid_control_slave_waits_for_read <= sysid_control_slave_in_a_read_cycle AND sysid_control_slave_begins_xfer;
  --sysid_control_slave_in_a_read_cycle assignment, which is an e_assign
  sysid_control_slave_in_a_read_cycle <= internal_peripheral_bridge_m1_granted_sysid_control_slave AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sysid_control_slave_in_a_read_cycle;
  --sysid_control_slave_waits_for_write in a cycle, which is an e_mux
  sysid_control_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysid_control_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sysid_control_slave_in_a_write_cycle assignment, which is an e_assign
  sysid_control_slave_in_a_write_cycle <= internal_peripheral_bridge_m1_granted_sysid_control_slave AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sysid_control_slave_in_a_write_cycle;
  wait_for_sysid_control_slave_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  peripheral_bridge_m1_granted_sysid_control_slave <= internal_peripheral_bridge_m1_granted_sysid_control_slave;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_qualified_request_sysid_control_slave <= internal_peripheral_bridge_m1_qualified_request_sysid_control_slave;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_requests_sysid_control_slave <= internal_peripheral_bridge_m1_requests_sysid_control_slave;
--synthesis translate_off
    --sysid/control_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --peripheral_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line118 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_peripheral_bridge_m1_requests_sysid_control_slave AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line118, now);
          write(write_line118, string'(": "));
          write(write_line118, string'("peripheral_bridge/m1 drove 0 on its 'burstcount' port while accessing slave sysid/control_slave"));
          write(output, write_line118.all);
          deallocate (write_line118);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity systimer_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                 signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                 signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read : IN STD_LOGIC;
                 signal peripheral_bridge_m1_write : IN STD_LOGIC;
                 signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal systimer_s1_irq : IN STD_LOGIC;
                 signal systimer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal d1_systimer_s1_end_xfer : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_granted_systimer_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_systimer_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_systimer_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_requests_systimer_s1 : OUT STD_LOGIC;
                 signal systimer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal systimer_s1_chipselect : OUT STD_LOGIC;
                 signal systimer_s1_irq_from_sa : OUT STD_LOGIC;
                 signal systimer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal systimer_s1_reset_n : OUT STD_LOGIC;
                 signal systimer_s1_write_n : OUT STD_LOGIC;
                 signal systimer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity systimer_s1_arbitrator;


architecture europa of systimer_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_systimer_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_granted_systimer_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_qualified_request_systimer_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_requests_systimer_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal peripheral_bridge_m1_continuerequest :  STD_LOGIC;
                signal peripheral_bridge_m1_saved_grant_systimer_s1 :  STD_LOGIC;
                signal shifted_address_to_systimer_s1_from_peripheral_bridge_m1 :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal systimer_s1_allgrants :  STD_LOGIC;
                signal systimer_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal systimer_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal systimer_s1_any_continuerequest :  STD_LOGIC;
                signal systimer_s1_arb_counter_enable :  STD_LOGIC;
                signal systimer_s1_arb_share_counter :  STD_LOGIC;
                signal systimer_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal systimer_s1_arb_share_set_values :  STD_LOGIC;
                signal systimer_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal systimer_s1_begins_xfer :  STD_LOGIC;
                signal systimer_s1_end_xfer :  STD_LOGIC;
                signal systimer_s1_firsttransfer :  STD_LOGIC;
                signal systimer_s1_grant_vector :  STD_LOGIC;
                signal systimer_s1_in_a_read_cycle :  STD_LOGIC;
                signal systimer_s1_in_a_write_cycle :  STD_LOGIC;
                signal systimer_s1_master_qreq_vector :  STD_LOGIC;
                signal systimer_s1_non_bursting_master_requests :  STD_LOGIC;
                signal systimer_s1_reg_firsttransfer :  STD_LOGIC;
                signal systimer_s1_slavearbiterlockenable :  STD_LOGIC;
                signal systimer_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal systimer_s1_unreg_firsttransfer :  STD_LOGIC;
                signal systimer_s1_waits_for_read :  STD_LOGIC;
                signal systimer_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_systimer_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT systimer_s1_end_xfer;
    end if;

  end process;

  systimer_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_peripheral_bridge_m1_qualified_request_systimer_s1);
  --assign systimer_s1_readdata_from_sa = systimer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  systimer_s1_readdata_from_sa <= systimer_s1_readdata;
  internal_peripheral_bridge_m1_requests_systimer_s1 <= to_std_logic(((Std_Logic_Vector'(peripheral_bridge_m1_address_to_slave(12 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("0000000100000")))) AND peripheral_bridge_m1_chipselect;
  --systimer_s1_arb_share_counter set values, which is an e_mux
  systimer_s1_arb_share_set_values <= std_logic'('1');
  --systimer_s1_non_bursting_master_requests mux, which is an e_mux
  systimer_s1_non_bursting_master_requests <= internal_peripheral_bridge_m1_requests_systimer_s1;
  --systimer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  systimer_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --systimer_s1_arb_share_counter_next_value assignment, which is an e_assign
  systimer_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(systimer_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(systimer_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(systimer_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(systimer_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --systimer_s1_allgrants all slave grants, which is an e_mux
  systimer_s1_allgrants <= systimer_s1_grant_vector;
  --systimer_s1_end_xfer assignment, which is an e_assign
  systimer_s1_end_xfer <= NOT ((systimer_s1_waits_for_read OR systimer_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_systimer_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_systimer_s1 <= systimer_s1_end_xfer AND (((NOT systimer_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --systimer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  systimer_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_systimer_s1 AND systimer_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_systimer_s1 AND NOT systimer_s1_non_bursting_master_requests));
  --systimer_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      systimer_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(systimer_s1_arb_counter_enable) = '1' then 
        systimer_s1_arb_share_counter <= systimer_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --systimer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      systimer_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((systimer_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_systimer_s1)) OR ((end_xfer_arb_share_counter_term_systimer_s1 AND NOT systimer_s1_non_bursting_master_requests)))) = '1' then 
        systimer_s1_slavearbiterlockenable <= systimer_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --peripheral_bridge/m1 systimer/s1 arbiterlock, which is an e_assign
  peripheral_bridge_m1_arbiterlock <= systimer_s1_slavearbiterlockenable AND peripheral_bridge_m1_continuerequest;
  --systimer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  systimer_s1_slavearbiterlockenable2 <= systimer_s1_arb_share_counter_next_value;
  --peripheral_bridge/m1 systimer/s1 arbiterlock2, which is an e_assign
  peripheral_bridge_m1_arbiterlock2 <= systimer_s1_slavearbiterlockenable2 AND peripheral_bridge_m1_continuerequest;
  --systimer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  systimer_s1_any_continuerequest <= std_logic'('1');
  --peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  peripheral_bridge_m1_continuerequest <= std_logic'('1');
  internal_peripheral_bridge_m1_qualified_request_systimer_s1 <= internal_peripheral_bridge_m1_requests_systimer_s1 AND NOT ((((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid peripheral_bridge_m1_read_data_valid_systimer_s1, which is an e_mux
  peripheral_bridge_m1_read_data_valid_systimer_s1 <= (internal_peripheral_bridge_m1_granted_systimer_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect))) AND NOT systimer_s1_waits_for_read;
  --systimer_s1_writedata mux, which is an e_mux
  systimer_s1_writedata <= peripheral_bridge_m1_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_peripheral_bridge_m1_granted_systimer_s1 <= internal_peripheral_bridge_m1_qualified_request_systimer_s1;
  --peripheral_bridge/m1 saved-grant systimer/s1, which is an e_assign
  peripheral_bridge_m1_saved_grant_systimer_s1 <= internal_peripheral_bridge_m1_requests_systimer_s1;
  --allow new arb cycle for systimer/s1, which is an e_assign
  systimer_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  systimer_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  systimer_s1_master_qreq_vector <= std_logic'('1');
  --systimer_s1_reset_n assignment, which is an e_assign
  systimer_s1_reset_n <= reset_n;
  systimer_s1_chipselect <= internal_peripheral_bridge_m1_granted_systimer_s1;
  --systimer_s1_firsttransfer first transaction, which is an e_assign
  systimer_s1_firsttransfer <= A_WE_StdLogic((std_logic'(systimer_s1_begins_xfer) = '1'), systimer_s1_unreg_firsttransfer, systimer_s1_reg_firsttransfer);
  --systimer_s1_unreg_firsttransfer first transaction, which is an e_assign
  systimer_s1_unreg_firsttransfer <= NOT ((systimer_s1_slavearbiterlockenable AND systimer_s1_any_continuerequest));
  --systimer_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      systimer_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(systimer_s1_begins_xfer) = '1' then 
        systimer_s1_reg_firsttransfer <= systimer_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --systimer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  systimer_s1_beginbursttransfer_internal <= systimer_s1_begins_xfer;
  --~systimer_s1_write_n assignment, which is an e_mux
  systimer_s1_write_n <= NOT ((internal_peripheral_bridge_m1_granted_systimer_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect))));
  shifted_address_to_systimer_s1_from_peripheral_bridge_m1 <= peripheral_bridge_m1_address_to_slave;
  --systimer_s1_address mux, which is an e_mux
  systimer_s1_address <= A_EXT (A_SRL(shifted_address_to_systimer_s1_from_peripheral_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 3);
  --d1_systimer_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_systimer_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_systimer_s1_end_xfer <= systimer_s1_end_xfer;
    end if;

  end process;

  --systimer_s1_waits_for_read in a cycle, which is an e_mux
  systimer_s1_waits_for_read <= systimer_s1_in_a_read_cycle AND systimer_s1_begins_xfer;
  --systimer_s1_in_a_read_cycle assignment, which is an e_assign
  systimer_s1_in_a_read_cycle <= internal_peripheral_bridge_m1_granted_systimer_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= systimer_s1_in_a_read_cycle;
  --systimer_s1_waits_for_write in a cycle, which is an e_mux
  systimer_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(systimer_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --systimer_s1_in_a_write_cycle assignment, which is an e_assign
  systimer_s1_in_a_write_cycle <= internal_peripheral_bridge_m1_granted_systimer_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= systimer_s1_in_a_write_cycle;
  wait_for_systimer_s1_counter <= std_logic'('0');
  --assign systimer_s1_irq_from_sa = systimer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  systimer_s1_irq_from_sa <= systimer_s1_irq;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_granted_systimer_s1 <= internal_peripheral_bridge_m1_granted_systimer_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_qualified_request_systimer_s1 <= internal_peripheral_bridge_m1_qualified_request_systimer_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_requests_systimer_s1 <= internal_peripheral_bridge_m1_requests_systimer_s1;
--synthesis translate_off
    --systimer/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --peripheral_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line119 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_peripheral_bridge_m1_requests_systimer_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line119, now);
          write(write_line119, string'(": "));
          write(write_line119, string'("peripheral_bridge/m1 drove 0 on its 'burstcount' port while accessing slave systimer/s1"));
          write(output, write_line119.all);
          deallocate (write_line119);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sysuart_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                 signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                 signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read : IN STD_LOGIC;
                 signal peripheral_bridge_m1_write : IN STD_LOGIC;
                 signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sysuart_s1_dataavailable : IN STD_LOGIC;
                 signal sysuart_s1_irq : IN STD_LOGIC;
                 signal sysuart_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sysuart_s1_readyfordata : IN STD_LOGIC;

              -- outputs:
                 signal d1_sysuart_s1_end_xfer : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_granted_sysuart_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_sysuart_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_sysuart_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_requests_sysuart_s1 : OUT STD_LOGIC;
                 signal sysuart_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal sysuart_s1_begintransfer : OUT STD_LOGIC;
                 signal sysuart_s1_chipselect : OUT STD_LOGIC;
                 signal sysuart_s1_dataavailable_from_sa : OUT STD_LOGIC;
                 signal sysuart_s1_irq_from_sa : OUT STD_LOGIC;
                 signal sysuart_s1_read_n : OUT STD_LOGIC;
                 signal sysuart_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sysuart_s1_readyfordata_from_sa : OUT STD_LOGIC;
                 signal sysuart_s1_reset_n : OUT STD_LOGIC;
                 signal sysuart_s1_write_n : OUT STD_LOGIC;
                 signal sysuart_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity sysuart_s1_arbitrator;


architecture europa of sysuart_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sysuart_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_granted_sysuart_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_qualified_request_sysuart_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_requests_sysuart_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal peripheral_bridge_m1_continuerequest :  STD_LOGIC;
                signal peripheral_bridge_m1_saved_grant_sysuart_s1 :  STD_LOGIC;
                signal shifted_address_to_sysuart_s1_from_peripheral_bridge_m1 :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal sysuart_s1_allgrants :  STD_LOGIC;
                signal sysuart_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal sysuart_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sysuart_s1_any_continuerequest :  STD_LOGIC;
                signal sysuart_s1_arb_counter_enable :  STD_LOGIC;
                signal sysuart_s1_arb_share_counter :  STD_LOGIC;
                signal sysuart_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal sysuart_s1_arb_share_set_values :  STD_LOGIC;
                signal sysuart_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal sysuart_s1_begins_xfer :  STD_LOGIC;
                signal sysuart_s1_end_xfer :  STD_LOGIC;
                signal sysuart_s1_firsttransfer :  STD_LOGIC;
                signal sysuart_s1_grant_vector :  STD_LOGIC;
                signal sysuart_s1_in_a_read_cycle :  STD_LOGIC;
                signal sysuart_s1_in_a_write_cycle :  STD_LOGIC;
                signal sysuart_s1_master_qreq_vector :  STD_LOGIC;
                signal sysuart_s1_non_bursting_master_requests :  STD_LOGIC;
                signal sysuart_s1_reg_firsttransfer :  STD_LOGIC;
                signal sysuart_s1_slavearbiterlockenable :  STD_LOGIC;
                signal sysuart_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal sysuart_s1_unreg_firsttransfer :  STD_LOGIC;
                signal sysuart_s1_waits_for_read :  STD_LOGIC;
                signal sysuart_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_sysuart_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sysuart_s1_end_xfer;
    end if;

  end process;

  sysuart_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_peripheral_bridge_m1_qualified_request_sysuart_s1);
  --assign sysuart_s1_readdata_from_sa = sysuart_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sysuart_s1_readdata_from_sa <= sysuart_s1_readdata;
  internal_peripheral_bridge_m1_requests_sysuart_s1 <= to_std_logic(((Std_Logic_Vector'(peripheral_bridge_m1_address_to_slave(12 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("0000001000000")))) AND peripheral_bridge_m1_chipselect;
  --assign sysuart_s1_dataavailable_from_sa = sysuart_s1_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  sysuart_s1_dataavailable_from_sa <= sysuart_s1_dataavailable;
  --assign sysuart_s1_readyfordata_from_sa = sysuart_s1_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sysuart_s1_readyfordata_from_sa <= sysuart_s1_readyfordata;
  --sysuart_s1_arb_share_counter set values, which is an e_mux
  sysuart_s1_arb_share_set_values <= std_logic'('1');
  --sysuart_s1_non_bursting_master_requests mux, which is an e_mux
  sysuart_s1_non_bursting_master_requests <= internal_peripheral_bridge_m1_requests_sysuart_s1;
  --sysuart_s1_any_bursting_master_saved_grant mux, which is an e_mux
  sysuart_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --sysuart_s1_arb_share_counter_next_value assignment, which is an e_assign
  sysuart_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sysuart_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysuart_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(sysuart_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysuart_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --sysuart_s1_allgrants all slave grants, which is an e_mux
  sysuart_s1_allgrants <= sysuart_s1_grant_vector;
  --sysuart_s1_end_xfer assignment, which is an e_assign
  sysuart_s1_end_xfer <= NOT ((sysuart_s1_waits_for_read OR sysuart_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_sysuart_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sysuart_s1 <= sysuart_s1_end_xfer AND (((NOT sysuart_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sysuart_s1_arb_share_counter arbitration counter enable, which is an e_assign
  sysuart_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sysuart_s1 AND sysuart_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_sysuart_s1 AND NOT sysuart_s1_non_bursting_master_requests));
  --sysuart_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysuart_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(sysuart_s1_arb_counter_enable) = '1' then 
        sysuart_s1_arb_share_counter <= sysuart_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sysuart_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysuart_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sysuart_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_sysuart_s1)) OR ((end_xfer_arb_share_counter_term_sysuart_s1 AND NOT sysuart_s1_non_bursting_master_requests)))) = '1' then 
        sysuart_s1_slavearbiterlockenable <= sysuart_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --peripheral_bridge/m1 sysuart/s1 arbiterlock, which is an e_assign
  peripheral_bridge_m1_arbiterlock <= sysuart_s1_slavearbiterlockenable AND peripheral_bridge_m1_continuerequest;
  --sysuart_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sysuart_s1_slavearbiterlockenable2 <= sysuart_s1_arb_share_counter_next_value;
  --peripheral_bridge/m1 sysuart/s1 arbiterlock2, which is an e_assign
  peripheral_bridge_m1_arbiterlock2 <= sysuart_s1_slavearbiterlockenable2 AND peripheral_bridge_m1_continuerequest;
  --sysuart_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  sysuart_s1_any_continuerequest <= std_logic'('1');
  --peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  peripheral_bridge_m1_continuerequest <= std_logic'('1');
  internal_peripheral_bridge_m1_qualified_request_sysuart_s1 <= internal_peripheral_bridge_m1_requests_sysuart_s1 AND NOT ((((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid peripheral_bridge_m1_read_data_valid_sysuart_s1, which is an e_mux
  peripheral_bridge_m1_read_data_valid_sysuart_s1 <= (internal_peripheral_bridge_m1_granted_sysuart_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect))) AND NOT sysuart_s1_waits_for_read;
  --sysuart_s1_writedata mux, which is an e_mux
  sysuart_s1_writedata <= peripheral_bridge_m1_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_peripheral_bridge_m1_granted_sysuart_s1 <= internal_peripheral_bridge_m1_qualified_request_sysuart_s1;
  --peripheral_bridge/m1 saved-grant sysuart/s1, which is an e_assign
  peripheral_bridge_m1_saved_grant_sysuart_s1 <= internal_peripheral_bridge_m1_requests_sysuart_s1;
  --allow new arb cycle for sysuart/s1, which is an e_assign
  sysuart_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sysuart_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sysuart_s1_master_qreq_vector <= std_logic'('1');
  sysuart_s1_begintransfer <= sysuart_s1_begins_xfer;
  --sysuart_s1_reset_n assignment, which is an e_assign
  sysuart_s1_reset_n <= reset_n;
  sysuart_s1_chipselect <= internal_peripheral_bridge_m1_granted_sysuart_s1;
  --sysuart_s1_firsttransfer first transaction, which is an e_assign
  sysuart_s1_firsttransfer <= A_WE_StdLogic((std_logic'(sysuart_s1_begins_xfer) = '1'), sysuart_s1_unreg_firsttransfer, sysuart_s1_reg_firsttransfer);
  --sysuart_s1_unreg_firsttransfer first transaction, which is an e_assign
  sysuart_s1_unreg_firsttransfer <= NOT ((sysuart_s1_slavearbiterlockenable AND sysuart_s1_any_continuerequest));
  --sysuart_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysuart_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sysuart_s1_begins_xfer) = '1' then 
        sysuart_s1_reg_firsttransfer <= sysuart_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sysuart_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sysuart_s1_beginbursttransfer_internal <= sysuart_s1_begins_xfer;
  --~sysuart_s1_read_n assignment, which is an e_mux
  sysuart_s1_read_n <= NOT ((internal_peripheral_bridge_m1_granted_sysuart_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect))));
  --~sysuart_s1_write_n assignment, which is an e_mux
  sysuart_s1_write_n <= NOT ((internal_peripheral_bridge_m1_granted_sysuart_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect))));
  shifted_address_to_sysuart_s1_from_peripheral_bridge_m1 <= peripheral_bridge_m1_address_to_slave;
  --sysuart_s1_address mux, which is an e_mux
  sysuart_s1_address <= A_EXT (A_SRL(shifted_address_to_sysuart_s1_from_peripheral_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 3);
  --d1_sysuart_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sysuart_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sysuart_s1_end_xfer <= sysuart_s1_end_xfer;
    end if;

  end process;

  --sysuart_s1_waits_for_read in a cycle, which is an e_mux
  sysuart_s1_waits_for_read <= sysuart_s1_in_a_read_cycle AND sysuart_s1_begins_xfer;
  --sysuart_s1_in_a_read_cycle assignment, which is an e_assign
  sysuart_s1_in_a_read_cycle <= internal_peripheral_bridge_m1_granted_sysuart_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sysuart_s1_in_a_read_cycle;
  --sysuart_s1_waits_for_write in a cycle, which is an e_mux
  sysuart_s1_waits_for_write <= sysuart_s1_in_a_write_cycle AND sysuart_s1_begins_xfer;
  --sysuart_s1_in_a_write_cycle assignment, which is an e_assign
  sysuart_s1_in_a_write_cycle <= internal_peripheral_bridge_m1_granted_sysuart_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sysuart_s1_in_a_write_cycle;
  wait_for_sysuart_s1_counter <= std_logic'('0');
  --assign sysuart_s1_irq_from_sa = sysuart_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  sysuart_s1_irq_from_sa <= sysuart_s1_irq;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_granted_sysuart_s1 <= internal_peripheral_bridge_m1_granted_sysuart_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_qualified_request_sysuart_s1 <= internal_peripheral_bridge_m1_qualified_request_sysuart_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_requests_sysuart_s1 <= internal_peripheral_bridge_m1_requests_sysuart_s1;
--synthesis translate_off
    --sysuart/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --peripheral_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line120 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_peripheral_bridge_m1_requests_sysuart_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line120, now);
          write(write_line120, string'(": "));
          write(write_line120, string'("peripheral_bridge/m1 drove 0 on its 'burstcount' port while accessing slave sysuart/s1"));
          write(output, write_line120.all);
          deallocate (write_line120);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity vga_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                 signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                 signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal peripheral_bridge_m1_read : IN STD_LOGIC;
                 signal peripheral_bridge_m1_write : IN STD_LOGIC;
                 signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal vga_s1_irq : IN STD_LOGIC;
                 signal vga_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal d1_vga_s1_end_xfer : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_granted_vga_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_qualified_request_vga_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_read_data_valid_vga_s1 : OUT STD_LOGIC;
                 signal peripheral_bridge_m1_requests_vga_s1 : OUT STD_LOGIC;
                 signal vga_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal vga_s1_irq_from_sa : OUT STD_LOGIC;
                 signal vga_s1_read : OUT STD_LOGIC;
                 signal vga_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal vga_s1_write : OUT STD_LOGIC;
                 signal vga_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity vga_s1_arbitrator;


architecture europa of vga_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_vga_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_granted_vga_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_qualified_request_vga_s1 :  STD_LOGIC;
                signal internal_peripheral_bridge_m1_requests_vga_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock :  STD_LOGIC;
                signal peripheral_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal peripheral_bridge_m1_continuerequest :  STD_LOGIC;
                signal peripheral_bridge_m1_saved_grant_vga_s1 :  STD_LOGIC;
                signal shifted_address_to_vga_s1_from_peripheral_bridge_m1 :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal vga_s1_allgrants :  STD_LOGIC;
                signal vga_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal vga_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal vga_s1_any_continuerequest :  STD_LOGIC;
                signal vga_s1_arb_counter_enable :  STD_LOGIC;
                signal vga_s1_arb_share_counter :  STD_LOGIC;
                signal vga_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal vga_s1_arb_share_set_values :  STD_LOGIC;
                signal vga_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal vga_s1_begins_xfer :  STD_LOGIC;
                signal vga_s1_end_xfer :  STD_LOGIC;
                signal vga_s1_firsttransfer :  STD_LOGIC;
                signal vga_s1_grant_vector :  STD_LOGIC;
                signal vga_s1_in_a_read_cycle :  STD_LOGIC;
                signal vga_s1_in_a_write_cycle :  STD_LOGIC;
                signal vga_s1_master_qreq_vector :  STD_LOGIC;
                signal vga_s1_non_bursting_master_requests :  STD_LOGIC;
                signal vga_s1_reg_firsttransfer :  STD_LOGIC;
                signal vga_s1_slavearbiterlockenable :  STD_LOGIC;
                signal vga_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal vga_s1_unreg_firsttransfer :  STD_LOGIC;
                signal vga_s1_waits_for_read :  STD_LOGIC;
                signal vga_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_vga_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT vga_s1_end_xfer;
    end if;

  end process;

  vga_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_peripheral_bridge_m1_qualified_request_vga_s1);
  --assign vga_s1_readdata_from_sa = vga_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  vga_s1_readdata_from_sa <= vga_s1_readdata;
  internal_peripheral_bridge_m1_requests_vga_s1 <= to_std_logic(((Std_Logic_Vector'(peripheral_bridge_m1_address_to_slave(12 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("0100000000000")))) AND peripheral_bridge_m1_chipselect;
  --vga_s1_arb_share_counter set values, which is an e_mux
  vga_s1_arb_share_set_values <= std_logic'('1');
  --vga_s1_non_bursting_master_requests mux, which is an e_mux
  vga_s1_non_bursting_master_requests <= internal_peripheral_bridge_m1_requests_vga_s1;
  --vga_s1_any_bursting_master_saved_grant mux, which is an e_mux
  vga_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --vga_s1_arb_share_counter_next_value assignment, which is an e_assign
  vga_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(vga_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(vga_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(vga_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(vga_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --vga_s1_allgrants all slave grants, which is an e_mux
  vga_s1_allgrants <= vga_s1_grant_vector;
  --vga_s1_end_xfer assignment, which is an e_assign
  vga_s1_end_xfer <= NOT ((vga_s1_waits_for_read OR vga_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_vga_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_vga_s1 <= vga_s1_end_xfer AND (((NOT vga_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --vga_s1_arb_share_counter arbitration counter enable, which is an e_assign
  vga_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_vga_s1 AND vga_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_vga_s1 AND NOT vga_s1_non_bursting_master_requests));
  --vga_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      vga_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(vga_s1_arb_counter_enable) = '1' then 
        vga_s1_arb_share_counter <= vga_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --vga_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      vga_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((vga_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_vga_s1)) OR ((end_xfer_arb_share_counter_term_vga_s1 AND NOT vga_s1_non_bursting_master_requests)))) = '1' then 
        vga_s1_slavearbiterlockenable <= vga_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --peripheral_bridge/m1 vga/s1 arbiterlock, which is an e_assign
  peripheral_bridge_m1_arbiterlock <= vga_s1_slavearbiterlockenable AND peripheral_bridge_m1_continuerequest;
  --vga_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  vga_s1_slavearbiterlockenable2 <= vga_s1_arb_share_counter_next_value;
  --peripheral_bridge/m1 vga/s1 arbiterlock2, which is an e_assign
  peripheral_bridge_m1_arbiterlock2 <= vga_s1_slavearbiterlockenable2 AND peripheral_bridge_m1_continuerequest;
  --vga_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  vga_s1_any_continuerequest <= std_logic'('1');
  --peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  peripheral_bridge_m1_continuerequest <= std_logic'('1');
  internal_peripheral_bridge_m1_qualified_request_vga_s1 <= internal_peripheral_bridge_m1_requests_vga_s1 AND NOT ((((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid peripheral_bridge_m1_read_data_valid_vga_s1, which is an e_mux
  peripheral_bridge_m1_read_data_valid_vga_s1 <= (internal_peripheral_bridge_m1_granted_vga_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect))) AND NOT vga_s1_waits_for_read;
  --vga_s1_writedata mux, which is an e_mux
  vga_s1_writedata <= peripheral_bridge_m1_writedata;
  --master is always granted when requested
  internal_peripheral_bridge_m1_granted_vga_s1 <= internal_peripheral_bridge_m1_qualified_request_vga_s1;
  --peripheral_bridge/m1 saved-grant vga/s1, which is an e_assign
  peripheral_bridge_m1_saved_grant_vga_s1 <= internal_peripheral_bridge_m1_requests_vga_s1;
  --allow new arb cycle for vga/s1, which is an e_assign
  vga_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  vga_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  vga_s1_master_qreq_vector <= std_logic'('1');
  --vga_s1_firsttransfer first transaction, which is an e_assign
  vga_s1_firsttransfer <= A_WE_StdLogic((std_logic'(vga_s1_begins_xfer) = '1'), vga_s1_unreg_firsttransfer, vga_s1_reg_firsttransfer);
  --vga_s1_unreg_firsttransfer first transaction, which is an e_assign
  vga_s1_unreg_firsttransfer <= NOT ((vga_s1_slavearbiterlockenable AND vga_s1_any_continuerequest));
  --vga_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      vga_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(vga_s1_begins_xfer) = '1' then 
        vga_s1_reg_firsttransfer <= vga_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --vga_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  vga_s1_beginbursttransfer_internal <= vga_s1_begins_xfer;
  --vga_s1_read assignment, which is an e_mux
  vga_s1_read <= internal_peripheral_bridge_m1_granted_vga_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --vga_s1_write assignment, which is an e_mux
  vga_s1_write <= internal_peripheral_bridge_m1_granted_vga_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect));
  shifted_address_to_vga_s1_from_peripheral_bridge_m1 <= peripheral_bridge_m1_address_to_slave;
  --vga_s1_address mux, which is an e_mux
  vga_s1_address <= A_EXT (A_SRL(shifted_address_to_vga_s1_from_peripheral_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_vga_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_vga_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_vga_s1_end_xfer <= vga_s1_end_xfer;
    end if;

  end process;

  --vga_s1_waits_for_read in a cycle, which is an e_mux
  vga_s1_waits_for_read <= vga_s1_in_a_read_cycle AND vga_s1_begins_xfer;
  --vga_s1_in_a_read_cycle assignment, which is an e_assign
  vga_s1_in_a_read_cycle <= internal_peripheral_bridge_m1_granted_vga_s1 AND ((peripheral_bridge_m1_read AND peripheral_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= vga_s1_in_a_read_cycle;
  --vga_s1_waits_for_write in a cycle, which is an e_mux
  vga_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(vga_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --vga_s1_in_a_write_cycle assignment, which is an e_assign
  vga_s1_in_a_write_cycle <= internal_peripheral_bridge_m1_granted_vga_s1 AND ((peripheral_bridge_m1_write AND peripheral_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= vga_s1_in_a_write_cycle;
  wait_for_vga_s1_counter <= std_logic'('0');
  --assign vga_s1_irq_from_sa = vga_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  vga_s1_irq_from_sa <= vga_s1_irq;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_granted_vga_s1 <= internal_peripheral_bridge_m1_granted_vga_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_qualified_request_vga_s1 <= internal_peripheral_bridge_m1_qualified_request_vga_s1;
  --vhdl renameroo for output signals
  peripheral_bridge_m1_requests_vga_s1 <= internal_peripheral_bridge_m1_requests_vga_s1;
--synthesis translate_off
    --vga/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --peripheral_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line121 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_peripheral_bridge_m1_requests_vga_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(peripheral_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line121, now);
          write(write_line121, string'(": "));
          write(write_line121, string'("peripheral_bridge/m1 drove 0 on its 'burstcount' port while accessing slave vga/s1"));
          write(output, write_line121.all);
          deallocate (write_line121);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity vga_m1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_nios2_fpu_burst_0_upstream_end_xfer : IN STD_LOGIC;
                 signal nios2_fpu_burst_0_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal nios2_fpu_burst_0_upstream_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal vga_m1_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal vga_m1_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal vga_m1_granted_nios2_fpu_burst_0_upstream : IN STD_LOGIC;
                 signal vga_m1_qualified_request_nios2_fpu_burst_0_upstream : IN STD_LOGIC;
                 signal vga_m1_read : IN STD_LOGIC;
                 signal vga_m1_read_data_valid_nios2_fpu_burst_0_upstream : IN STD_LOGIC;
                 signal vga_m1_read_data_valid_nios2_fpu_burst_0_upstream_shift_register : IN STD_LOGIC;
                 signal vga_m1_requests_nios2_fpu_burst_0_upstream : IN STD_LOGIC;

              -- outputs:
                 signal vga_m1_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal vga_m1_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal vga_m1_latency_counter : OUT STD_LOGIC;
                 signal vga_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal vga_m1_readdatavalid : OUT STD_LOGIC;
                 signal vga_m1_reset : OUT STD_LOGIC;
                 signal vga_m1_waitrequest : OUT STD_LOGIC
              );
end entity vga_m1_arbitrator;


architecture europa of vga_m1_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dbs_rdv_count_enable :  STD_LOGIC;
                signal dbs_rdv_counter_overflow :  STD_LOGIC;
                signal internal_vga_m1_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_vga_m1_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_vga_m1_waitrequest :  STD_LOGIC;
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal pre_flush_vga_m1_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal vga_m1_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal vga_m1_burstcount_last_time :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal vga_m1_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal vga_m1_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal vga_m1_dbs_rdv_counter_inc :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal vga_m1_next_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal vga_m1_read_last_time :  STD_LOGIC;
                signal vga_m1_run :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((vga_m1_qualified_request_nios2_fpu_burst_0_upstream OR NOT vga_m1_requests_nios2_fpu_burst_0_upstream)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT vga_m1_qualified_request_nios2_fpu_burst_0_upstream OR NOT vga_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_0_upstream_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(vga_m1_read)))))))));
  --cascaded wait assignment, which is an e_assign
  vga_m1_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_vga_m1_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("0000000") & vga_m1_address(24 DOWNTO 0));
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_vga_m1_readdatavalid <= vga_m1_read_data_valid_nios2_fpu_burst_0_upstream AND dbs_rdv_counter_overflow;
  --latent slave read data valid which is not flushed, which is an e_mux
  vga_m1_readdatavalid <= Vector_To_Std_Logic((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_vga_m1_readdatavalid)))));
  --input to latent dbs-16 stored 0, which is an e_mux
  p1_dbs_latent_16_reg_segment_0 <= nios2_fpu_burst_0_upstream_readdata_from_sa;
  --dbs register for latent dbs-16 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_16_reg_segment_0 <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((vga_m1_dbs_rdv_counter(1))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
      end if;
    end if;

  end process;

  --vga/m1 readdata mux, which is an e_mux
  vga_m1_readdata <= Std_Logic_Vector'(nios2_fpu_burst_0_upstream_readdata_from_sa(15 DOWNTO 0) & dbs_latent_16_reg_segment_0);
  --actual waitrequest port, which is an e_assign
  internal_vga_m1_waitrequest <= NOT vga_m1_run;
  --latent max counter, which is an e_assign
  vga_m1_latency_counter <= std_logic'('0');
  --~vga_m1_reset assignment, which is an e_assign
  vga_m1_reset <= NOT reset_n;
  --dbs count increment, which is an e_mux
  vga_m1_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((vga_m1_requests_nios2_fpu_burst_0_upstream)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000000")), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_vga_m1_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_vga_m1_dbs_address)) + (std_logic_vector'("0") & (vga_m1_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_vga_m1_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_vga_m1_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --p1 dbs rdv counter, which is an e_assign
  vga_m1_next_dbs_rdv_counter <= A_EXT (((std_logic_vector'("0") & (vga_m1_dbs_rdv_counter)) + (std_logic_vector'("0") & (vga_m1_dbs_rdv_counter_inc))), 2);
  --vga_m1_rdv_inc_mux, which is an e_mux
  vga_m1_dbs_rdv_counter_inc <= std_logic_vector'("10");
  --master any slave rdv, which is an e_mux
  dbs_rdv_count_enable <= vga_m1_read_data_valid_nios2_fpu_burst_0_upstream;
  --dbs rdv counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      vga_m1_dbs_rdv_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_rdv_count_enable) = '1' then 
        vga_m1_dbs_rdv_counter <= vga_m1_next_dbs_rdv_counter;
      end if;
    end if;

  end process;

  --dbs rdv counter overflow, which is an e_assign
  dbs_rdv_counter_overflow <= vga_m1_dbs_rdv_counter(1) AND NOT vga_m1_next_dbs_rdv_counter(1);
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic(((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((vga_m1_granted_nios2_fpu_burst_0_upstream AND vga_m1_read)))) AND std_logic_vector'("00000000000000000000000000000000")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT nios2_fpu_burst_0_upstream_waitrequest_from_sa)))));
  --vhdl renameroo for output signals
  vga_m1_address_to_slave <= internal_vga_m1_address_to_slave;
  --vhdl renameroo for output signals
  vga_m1_dbs_address <= internal_vga_m1_dbs_address;
  --vhdl renameroo for output signals
  vga_m1_waitrequest <= internal_vga_m1_waitrequest;
--synthesis translate_off
    --vga_m1_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        vga_m1_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        vga_m1_address_last_time <= vga_m1_address;
      end if;

    end process;

    --vga/m1 waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_vga_m1_waitrequest AND (vga_m1_read);
      end if;

    end process;

    --vga_m1_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line122 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((vga_m1_address /= vga_m1_address_last_time))))) = '1' then 
          write(write_line122, now);
          write(write_line122, string'(": "));
          write(write_line122, string'("vga_m1_address did not heed wait!!!"));
          write(output, write_line122.all);
          deallocate (write_line122);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --vga_m1_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        vga_m1_burstcount_last_time <= std_logic_vector'("0000000000");
      elsif clk'event and clk = '1' then
        vga_m1_burstcount_last_time <= vga_m1_burstcount;
      end if;

    end process;

    --vga_m1_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line123 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((vga_m1_burstcount /= vga_m1_burstcount_last_time))))) = '1' then 
          write(write_line123, now);
          write(write_line123, string'(": "));
          write(write_line123, string'("vga_m1_burstcount did not heed wait!!!"));
          write(output, write_line123.all);
          deallocate (write_line123);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --vga_m1_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        vga_m1_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        vga_m1_read_last_time <= vga_m1_read;
      end if;

    end process;

    --vga_m1_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line124 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(vga_m1_read) /= std_logic'(vga_m1_read_last_time)))))) = '1' then 
          write(write_line124, now);
          write(write_line124, string'(": "));
          write(write_line124, string'("vga_m1_read did not heed wait!!!"));
          write(output, write_line124.all);
          deallocate (write_line124);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_fpu_reset_peri_clk_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity nios2_fpu_reset_peri_clk_domain_synch_module;


architecture europa of nios2_fpu_reset_peri_clk_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_fpu_reset_core_clk_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity nios2_fpu_reset_core_clk_domain_synch_module;


architecture europa of nios2_fpu_reset_core_clk_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity nios2_fpu is 
        port (
              -- 1) global signals:
                 signal core_clk : IN STD_LOGIC;
                 signal peri_clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- the_dipsw
                 signal in_port_to_the_dipsw : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

              -- the_gpio0
                 signal bidir_port_to_and_from_the_gpio0 : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- the_led
                 signal out_port_from_the_led : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_mmcdma
                 signal MMC_CD_to_the_mmcdma : IN STD_LOGIC;
                 signal MMC_SCK_from_the_mmcdma : OUT STD_LOGIC;
                 signal MMC_SDI_to_the_mmcdma : IN STD_LOGIC;
                 signal MMC_SDO_from_the_mmcdma : OUT STD_LOGIC;
                 signal MMC_WP_to_the_mmcdma : IN STD_LOGIC;
                 signal MMC_nCS_from_the_mmcdma : OUT STD_LOGIC;

              -- the_psw
                 signal in_port_to_the_psw : IN STD_LOGIC_VECTOR (1 DOWNTO 0);

              -- the_sdram
                 signal zs_addr_from_the_sdram : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal zs_ba_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal zs_cas_n_from_the_sdram : OUT STD_LOGIC;
                 signal zs_cke_from_the_sdram : OUT STD_LOGIC;
                 signal zs_cs_n_from_the_sdram : OUT STD_LOGIC;
                 signal zs_dq_to_and_from_the_sdram : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal zs_dqm_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal zs_ras_n_from_the_sdram : OUT STD_LOGIC;
                 signal zs_we_n_from_the_sdram : OUT STD_LOGIC;

              -- the_spu
                 signal AUD_L_from_the_spu : OUT STD_LOGIC;
                 signal AUD_R_from_the_spu : OUT STD_LOGIC;
                 signal DAC_BCLK_from_the_spu : OUT STD_LOGIC;
                 signal DAC_DATA_from_the_spu : OUT STD_LOGIC;
                 signal DAC_LRCK_from_the_spu : OUT STD_LOGIC;
                 signal SPDIF_from_the_spu : OUT STD_LOGIC;
                 signal clk_128fs_to_the_spu : IN STD_LOGIC;

              -- the_sysuart
                 signal rxd_to_the_sysuart : IN STD_LOGIC;
                 signal txd_from_the_sysuart : OUT STD_LOGIC;

              -- the_vga
                 signal video_bout_from_the_vga : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal video_clk_to_the_vga : IN STD_LOGIC;
                 signal video_enable_from_the_vga : OUT STD_LOGIC;
                 signal video_gout_from_the_vga : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal video_hsync_n_from_the_vga : OUT STD_LOGIC;
                 signal video_rout_from_the_vga : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal video_vsync_n_from_the_vga : OUT STD_LOGIC
              );
end entity nios2_fpu;


architecture europa of nios2_fpu is
component dipsw_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal dipsw_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                    signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                    signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read : IN STD_LOGIC;
                    signal peripheral_bridge_m1_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_dipsw_s1_end_xfer : OUT STD_LOGIC;
                    signal dipsw_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal dipsw_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal dipsw_s1_reset_n : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_granted_dipsw_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_dipsw_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_dipsw_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_requests_dipsw_s1 : OUT STD_LOGIC
                 );
end component dipsw_s1_arbitrator;

component dipsw is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal in_port : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component dipsw;

component gpio0_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal gpio0_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                    signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                    signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read : IN STD_LOGIC;
                    signal peripheral_bridge_m1_write : IN STD_LOGIC;
                    signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_gpio0_s1_end_xfer : OUT STD_LOGIC;
                    signal gpio0_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal gpio0_s1_chipselect : OUT STD_LOGIC;
                    signal gpio0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal gpio0_s1_reset_n : OUT STD_LOGIC;
                    signal gpio0_s1_write_n : OUT STD_LOGIC;
                    signal gpio0_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal peripheral_bridge_m1_granted_gpio0_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_gpio0_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_gpio0_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_requests_gpio0_s1 : OUT STD_LOGIC
                 );
end component gpio0_s1_arbitrator;

component gpio0 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal bidir_port : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component gpio0;

component ipl_memory_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal ipl_memory_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_6_downstream_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_burst_6_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_6_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_6_downstream_latency_counter : IN STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_7_downstream_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_burst_7_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_7_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_7_downstream_latency_counter : IN STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_ipl_memory_s1_end_xfer : OUT STD_LOGIC;
                    signal ipl_memory_s1_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal ipl_memory_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal ipl_memory_s1_chipselect : OUT STD_LOGIC;
                    signal ipl_memory_s1_clken : OUT STD_LOGIC;
                    signal ipl_memory_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ipl_memory_s1_reset : OUT STD_LOGIC;
                    signal ipl_memory_s1_write : OUT STD_LOGIC;
                    signal ipl_memory_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_requests_ipl_memory_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_granted_ipl_memory_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_requests_ipl_memory_s1 : OUT STD_LOGIC
                 );
end component ipl_memory_s1_arbitrator;

component ipl_memory is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal clken : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component ipl_memory;

component jtag_uart_avalon_jtag_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                    signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                    signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                    signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read : IN STD_LOGIC;
                    signal peripheral_bridge_m1_write : IN STD_LOGIC;
                    signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_jtag_uart_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_address : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC
                 );
end component jtag_uart_avalon_jtag_slave_arbitrator;

component jtag_uart is 
           port (
                 -- inputs:
                    signal av_address : IN STD_LOGIC;
                    signal av_chipselect : IN STD_LOGIC;
                    signal av_read_n : IN STD_LOGIC;
                    signal av_write_n : IN STD_LOGIC;
                    signal av_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal rst_n : IN STD_LOGIC;

                 -- outputs:
                    signal av_irq : OUT STD_LOGIC;
                    signal av_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal av_waitrequest : OUT STD_LOGIC;
                    signal dataavailable : OUT STD_LOGIC;
                    signal readyfordata : OUT STD_LOGIC
                 );
end component jtag_uart;

component led_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal led_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                    signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                    signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read : IN STD_LOGIC;
                    signal peripheral_bridge_m1_write : IN STD_LOGIC;
                    signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_led_s1_end_xfer : OUT STD_LOGIC;
                    signal led_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal led_s1_chipselect : OUT STD_LOGIC;
                    signal led_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal led_s1_reset_n : OUT STD_LOGIC;
                    signal led_s1_write_n : OUT STD_LOGIC;
                    signal led_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal peripheral_bridge_m1_granted_led_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_led_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_led_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_requests_led_s1 : OUT STD_LOGIC
                 );
end component led_s1_arbitrator;

component led is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component led;

component mmcdma_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal mmcdma_s1_irq : IN STD_LOGIC;
                    signal mmcdma_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                    signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                    signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read : IN STD_LOGIC;
                    signal peripheral_bridge_m1_write : IN STD_LOGIC;
                    signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_mmcdma_s1_end_xfer : OUT STD_LOGIC;
                    signal mmcdma_s1_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal mmcdma_s1_chipselect : OUT STD_LOGIC;
                    signal mmcdma_s1_irq_from_sa : OUT STD_LOGIC;
                    signal mmcdma_s1_read : OUT STD_LOGIC;
                    signal mmcdma_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal mmcdma_s1_reset : OUT STD_LOGIC;
                    signal mmcdma_s1_wait_counter_eq_0 : OUT STD_LOGIC;
                    signal mmcdma_s1_write : OUT STD_LOGIC;
                    signal mmcdma_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal peripheral_bridge_m1_granted_mmcdma_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_mmcdma_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_mmcdma_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_requests_mmcdma_s1 : OUT STD_LOGIC
                 );
end component mmcdma_s1_arbitrator;

component mmcdma is 
           port (
                 -- inputs:
                    signal MMC_CD : IN STD_LOGIC;
                    signal MMC_SDI : IN STD_LOGIC;
                    signal MMC_WP : IN STD_LOGIC;
                    signal address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal MMC_SCK : OUT STD_LOGIC;
                    signal MMC_SDO : OUT STD_LOGIC;
                    signal MMC_nCS : OUT STD_LOGIC;
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component mmcdma;

component nios2_fast_fpu_jtag_debug_module_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fast_fpu_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_jtag_debug_module_resetrequest : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_address_to_slave : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal nios2_fpu_burst_4_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_4_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_4_downstream_debugaccess : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_latency_counter : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_5_downstream_address_to_slave : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal nios2_fpu_burst_5_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_5_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_5_downstream_debugaccess : IN STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_latency_counter : IN STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_nios2_fast_fpu_jtag_debug_module_end_xfer : OUT STD_LOGIC;
                    signal nios2_fast_fpu_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal nios2_fast_fpu_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                    signal nios2_fast_fpu_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fast_fpu_jtag_debug_module_chipselect : OUT STD_LOGIC;
                    signal nios2_fast_fpu_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                    signal nios2_fast_fpu_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_fast_fpu_jtag_debug_module_write : OUT STD_LOGIC;
                    signal nios2_fast_fpu_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module : OUT STD_LOGIC
                 );
end component nios2_fast_fpu_jtag_debug_module_arbitrator;

component nios2_fast_fpu_custom_instruction_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fast_fpu_custom_instruction_master_multi_n : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_fast_fpu_custom_instruction_master_multi_start : IN STD_LOGIC;
                    signal nios2_fast_fpu_fpoint_s1_done_from_sa : IN STD_LOGIC;
                    signal nios2_fast_fpu_fpoint_s1_result_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done_from_sa : IN STD_LOGIC;
                    signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_fast_fpu_custom_instruction_master_multi_done : OUT STD_LOGIC;
                    signal nios2_fast_fpu_custom_instruction_master_multi_result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_custom_instruction_master_reset_n : OUT STD_LOGIC;
                    signal nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_fpoint_s1 : OUT STD_LOGIC;
                    signal nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0 : OUT STD_LOGIC;
                    signal nios2_fast_fpu_fpoint_s1_select : OUT STD_LOGIC;
                    signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select : OUT STD_LOGIC
                 );
end component nios2_fast_fpu_custom_instruction_master_arbitrator;

component nios2_fast_fpu_data_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal core_clk : IN STD_LOGIC;
                    signal core_clk_reset_n : IN STD_LOGIC;
                    signal d1_nios2_fpu_burst_2_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_fpu_burst_5_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_fpu_burst_6_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_fpu_burst_8_upstream_end_xfer : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                    signal mmcdma_s1_irq_from_sa : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_address : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_write : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_2_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_2_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_fpu_burst_5_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_5_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_fpu_burst_6_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_6_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_fpu_burst_8_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_8_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal psw_s1_irq_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal spu_s1_irq_from_sa : IN STD_LOGIC;
                    signal systimer_s1_irq_from_sa : IN STD_LOGIC;
                    signal sysuart_s1_irq_from_sa : IN STD_LOGIC;
                    signal vga_s1_irq_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_fast_fpu_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_latency_counter : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_readdatavalid : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fast_fpu_data_master_arbitrator;

component nios2_fast_fpu_instruction_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_nios2_fpu_burst_1_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_fpu_burst_4_upstream_end_xfer : IN STD_LOGIC;
                    signal d1_nios2_fpu_burst_7_upstream_end_xfer : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_address : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal nios2_fast_fpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_1_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_4_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal nios2_fpu_burst_7_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_7_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_fast_fpu_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal nios2_fast_fpu_instruction_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fast_fpu_instruction_master_latency_counter : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_instruction_master_readdatavalid : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fast_fpu_instruction_master_arbitrator;

component nios2_fast_fpu is 
           port (
                 -- inputs:
                    signal A_ci_multi_done : IN STD_LOGIC;
                    signal A_ci_multi_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d_irq : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_readdatavalid : IN STD_LOGIC;
                    signal d_waitrequest : IN STD_LOGIC;
                    signal i_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_readdatavalid : IN STD_LOGIC;
                    signal i_waitrequest : IN STD_LOGIC;
                    signal jtag_debug_module_address : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal jtag_debug_module_begintransfer : IN STD_LOGIC;
                    signal jtag_debug_module_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal jtag_debug_module_debugaccess : IN STD_LOGIC;
                    signal jtag_debug_module_select : IN STD_LOGIC;
                    signal jtag_debug_module_write : IN STD_LOGIC;
                    signal jtag_debug_module_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal A_ci_multi_a : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal A_ci_multi_b : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal A_ci_multi_c : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal A_ci_multi_clk_en : OUT STD_LOGIC;
                    signal A_ci_multi_clock : OUT STD_LOGIC;
                    signal A_ci_multi_dataa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal A_ci_multi_datab : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal A_ci_multi_estatus : OUT STD_LOGIC;
                    signal A_ci_multi_ipending : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal A_ci_multi_n : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal A_ci_multi_readra : OUT STD_LOGIC;
                    signal A_ci_multi_readrb : OUT STD_LOGIC;
                    signal A_ci_multi_reset : OUT STD_LOGIC;
                    signal A_ci_multi_start : OUT STD_LOGIC;
                    signal A_ci_multi_status : OUT STD_LOGIC;
                    signal A_ci_multi_writerc : OUT STD_LOGIC;
                    signal d_address : OUT STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal d_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal d_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal d_read : OUT STD_LOGIC;
                    signal d_write : OUT STD_LOGIC;
                    signal d_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_address : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal i_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal i_read : OUT STD_LOGIC;
                    signal jtag_debug_module_debugaccess_to_roms : OUT STD_LOGIC;
                    signal jtag_debug_module_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_debug_module_resetrequest : OUT STD_LOGIC
                 );
end component nios2_fast_fpu;

component nios2_fast_fpu_fpoint_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fast_fpu_custom_instruction_master_multi_clk_en : IN STD_LOGIC;
                    signal nios2_fast_fpu_custom_instruction_master_multi_dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_custom_instruction_master_multi_datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_custom_instruction_master_multi_n : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_fpoint_s1 : IN STD_LOGIC;
                    signal nios2_fast_fpu_fpoint_s1_done : IN STD_LOGIC;
                    signal nios2_fast_fpu_fpoint_s1_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_fpoint_s1_select : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_fast_fpu_fpoint_s1_clk_en : OUT STD_LOGIC;
                    signal nios2_fast_fpu_fpoint_s1_dataa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_fpoint_s1_datab : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_fpoint_s1_done_from_sa : OUT STD_LOGIC;
                    signal nios2_fast_fpu_fpoint_s1_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fast_fpu_fpoint_s1_reset : OUT STD_LOGIC;
                    signal nios2_fast_fpu_fpoint_s1_result_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_fpoint_s1_start : OUT STD_LOGIC
                 );
end component nios2_fast_fpu_fpoint_s1_arbitrator;

component nios2_fast_fpu_fpoint is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clk_en : IN STD_LOGIC;
                    signal dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal n : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reset : IN STD_LOGIC;
                    signal start : IN STD_LOGIC;

                 -- outputs:
                    signal done : OUT STD_LOGIC;
                    signal result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component nios2_fast_fpu_fpoint;

component nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fast_fpu_custom_instruction_master_multi_clk_en : IN STD_LOGIC;
                    signal nios2_fast_fpu_custom_instruction_master_multi_dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_custom_instruction_master_multi_datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_custom_instruction_master_multi_n : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0 : IN STD_LOGIC;
                    signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done : IN STD_LOGIC;
                    signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_clk_en : OUT STD_LOGIC;
                    signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_dataa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_datab : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done_from_sa : OUT STD_LOGIC;
                    signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_n : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_reset : OUT STD_LOGIC;
                    signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_start : OUT STD_LOGIC
                 );
end component nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_arbitrator;

component nios2_fast_fpu_pixelsimd_inst is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clk_en : IN STD_LOGIC;
                    signal dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal n : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal reset : IN STD_LOGIC;
                    signal start : IN STD_LOGIC;

                 -- outputs:
                    signal done : OUT STD_LOGIC;
                    signal result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component nios2_fast_fpu_pixelsimd_inst;

component nios2_fpu_burst_0_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_0_upstream_readdatavalid : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal vga_m1_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal vga_m1_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal vga_m1_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal vga_m1_latency_counter : IN STD_LOGIC;
                    signal vga_m1_read : IN STD_LOGIC;

                 -- outputs:
                    signal d1_nios2_fpu_burst_0_upstream_end_xfer : OUT STD_LOGIC;
                    signal nios2_fpu_burst_0_upstream_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_0_upstream_burstcount : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal nios2_fpu_burst_0_upstream_byteaddress : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal nios2_fpu_burst_0_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fpu_burst_0_upstream_debugaccess : OUT STD_LOGIC;
                    signal nios2_fpu_burst_0_upstream_read : OUT STD_LOGIC;
                    signal nios2_fpu_burst_0_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_0_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_fpu_burst_0_upstream_write : OUT STD_LOGIC;
                    signal vga_m1_granted_nios2_fpu_burst_0_upstream : OUT STD_LOGIC;
                    signal vga_m1_qualified_request_nios2_fpu_burst_0_upstream : OUT STD_LOGIC;
                    signal vga_m1_read_data_valid_nios2_fpu_burst_0_upstream : OUT STD_LOGIC;
                    signal vga_m1_read_data_valid_nios2_fpu_burst_0_upstream_shift_register : OUT STD_LOGIC;
                    signal vga_m1_requests_nios2_fpu_burst_0_upstream : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_0_upstream_arbitrator;

component nios2_fpu_burst_0_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_0_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fpu_burst_0_downstream_granted_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_qualified_request_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_requests_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_fpu_burst_0_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_0_downstream_latency_counter : OUT STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_0_downstream_readdatavalid : OUT STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_reset_n : OUT STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_0_downstream_arbitrator;

component nios2_fpu_burst_0 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal downstream_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal downstream_burstcount : OUT STD_LOGIC;
                    signal downstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal downstream_debugaccess : OUT STD_LOGIC;
                    signal downstream_nativeaddress : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal downstream_read : OUT STD_LOGIC;
                    signal downstream_write : OUT STD_LOGIC;
                    signal downstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_0;

component nios2_fpu_burst_1_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal nios2_fast_fpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fast_fpu_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fast_fpu_instruction_master_latency_counter : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_1_upstream_readdatavalid : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_nios2_fpu_burst_1_upstream_end_xfer : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream : OUT STD_LOGIC;
                    signal nios2_fpu_burst_1_upstream_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_1_upstream_byteaddress : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal nios2_fpu_burst_1_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fpu_burst_1_upstream_debugaccess : OUT STD_LOGIC;
                    signal nios2_fpu_burst_1_upstream_read : OUT STD_LOGIC;
                    signal nios2_fpu_burst_1_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_1_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_fpu_burst_1_upstream_write : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_1_upstream_arbitrator;

component nios2_fpu_burst_1_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_1_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fpu_burst_1_downstream_granted_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_qualified_request_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_requests_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_fpu_burst_1_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_1_downstream_latency_counter : OUT STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_1_downstream_readdatavalid : OUT STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_reset_n : OUT STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_1_downstream_arbitrator;

component nios2_fpu_burst_1 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_1;

component nios2_fpu_burst_2_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_debugaccess : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_latency_counter : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_2_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_2_upstream_readdatavalid : IN STD_LOGIC;
                    signal nios2_fpu_burst_2_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_nios2_fpu_burst_2_upstream_end_xfer : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream : OUT STD_LOGIC;
                    signal nios2_fpu_burst_2_upstream_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_2_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_2_upstream_byteaddress : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal nios2_fpu_burst_2_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fpu_burst_2_upstream_debugaccess : OUT STD_LOGIC;
                    signal nios2_fpu_burst_2_upstream_read : OUT STD_LOGIC;
                    signal nios2_fpu_burst_2_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_2_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_fpu_burst_2_upstream_write : OUT STD_LOGIC;
                    signal nios2_fpu_burst_2_upstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component nios2_fpu_burst_2_upstream_arbitrator;

component nios2_fpu_burst_2_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_2_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fpu_burst_2_downstream_granted_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_qualified_request_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_requests_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_fpu_burst_2_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_2_downstream_latency_counter : OUT STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_2_downstream_readdatavalid : OUT STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_reset_n : OUT STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_2_downstream_arbitrator;

component nios2_fpu_burst_2 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_2;

component nios2_fpu_burst_3_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_upstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_3_upstream_readdatavalid : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal spu_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal spu_m1_burstcount : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal spu_m1_latency_counter : IN STD_LOGIC;
                    signal spu_m1_read : IN STD_LOGIC;

                 -- outputs:
                    signal d1_nios2_fpu_burst_3_upstream_end_xfer : OUT STD_LOGIC;
                    signal nios2_fpu_burst_3_upstream_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_3_upstream_burstcount : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_fpu_burst_3_upstream_byteaddress : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal nios2_fpu_burst_3_upstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fpu_burst_3_upstream_debugaccess : OUT STD_LOGIC;
                    signal nios2_fpu_burst_3_upstream_read : OUT STD_LOGIC;
                    signal nios2_fpu_burst_3_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_3_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_fpu_burst_3_upstream_write : OUT STD_LOGIC;
                    signal spu_m1_granted_nios2_fpu_burst_3_upstream : OUT STD_LOGIC;
                    signal spu_m1_qualified_request_nios2_fpu_burst_3_upstream : OUT STD_LOGIC;
                    signal spu_m1_read_data_valid_nios2_fpu_burst_3_upstream : OUT STD_LOGIC;
                    signal spu_m1_read_data_valid_nios2_fpu_burst_3_upstream_shift_register : OUT STD_LOGIC;
                    signal spu_m1_requests_nios2_fpu_burst_3_upstream : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_3_upstream_arbitrator;

component nios2_fpu_burst_3_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_3_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fpu_burst_3_downstream_granted_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_qualified_request_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_requests_sdram_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_fpu_burst_3_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_3_downstream_latency_counter : OUT STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_3_downstream_readdatavalid : OUT STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_reset_n : OUT STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_3_downstream_arbitrator;

component nios2_fpu_burst_3 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_3;

component nios2_fpu_burst_4_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal nios2_fast_fpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fast_fpu_instruction_master_latency_counter : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_4_upstream_readdatavalid : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_nios2_fpu_burst_4_upstream_end_xfer : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream : OUT STD_LOGIC;
                    signal nios2_fpu_burst_4_upstream_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal nios2_fpu_burst_4_upstream_byteaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_burst_4_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_4_upstream_debugaccess : OUT STD_LOGIC;
                    signal nios2_fpu_burst_4_upstream_read : OUT STD_LOGIC;
                    signal nios2_fpu_burst_4_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_4_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_fpu_burst_4_upstream_write : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_4_upstream_arbitrator;

component nios2_fpu_burst_4_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_nios2_fast_fpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal nios2_fast_fpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_4_downstream_address : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal nios2_fpu_burst_4_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_fpu_burst_4_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal nios2_fpu_burst_4_downstream_latency_counter : OUT STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_4_downstream_readdatavalid : OUT STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_reset_n : OUT STD_LOGIC;
                    signal nios2_fpu_burst_4_downstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_4_downstream_arbitrator;

component nios2_fpu_burst_4 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_4;

component nios2_fpu_burst_5_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_debugaccess : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_latency_counter : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_write : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_5_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_5_upstream_readdatavalid : IN STD_LOGIC;
                    signal nios2_fpu_burst_5_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_nios2_fpu_burst_5_upstream_end_xfer : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream : OUT STD_LOGIC;
                    signal nios2_fpu_burst_5_upstream_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal nios2_fpu_burst_5_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_5_upstream_byteaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_burst_5_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_5_upstream_debugaccess : OUT STD_LOGIC;
                    signal nios2_fpu_burst_5_upstream_read : OUT STD_LOGIC;
                    signal nios2_fpu_burst_5_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_5_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_fpu_burst_5_upstream_write : OUT STD_LOGIC;
                    signal nios2_fpu_burst_5_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component nios2_fpu_burst_5_upstream_arbitrator;

component nios2_fpu_burst_5_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_nios2_fast_fpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal nios2_fast_fpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_5_downstream_address : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal nios2_fpu_burst_5_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module : IN STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_fpu_burst_5_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal nios2_fpu_burst_5_downstream_latency_counter : OUT STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_5_downstream_readdatavalid : OUT STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_reset_n : OUT STD_LOGIC;
                    signal nios2_fpu_burst_5_downstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_5_downstream_arbitrator;

component nios2_fpu_burst_5 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_5;

component nios2_fpu_burst_6_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_debugaccess : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_latency_counter : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_write : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_6_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_6_upstream_readdatavalid : IN STD_LOGIC;
                    signal nios2_fpu_burst_6_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_nios2_fpu_burst_6_upstream_end_xfer : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream : OUT STD_LOGIC;
                    signal nios2_fpu_burst_6_upstream_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_burst_6_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_6_upstream_byteaddress : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal nios2_fpu_burst_6_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_6_upstream_debugaccess : OUT STD_LOGIC;
                    signal nios2_fpu_burst_6_upstream_read : OUT STD_LOGIC;
                    signal nios2_fpu_burst_6_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_6_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_fpu_burst_6_upstream_write : OUT STD_LOGIC;
                    signal nios2_fpu_burst_6_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component nios2_fpu_burst_6_upstream_arbitrator;

component nios2_fpu_burst_6_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_ipl_memory_s1_end_xfer : IN STD_LOGIC;
                    signal ipl_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_6_downstream_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_burst_6_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_requests_ipl_memory_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_fpu_burst_6_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_burst_6_downstream_latency_counter : OUT STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_6_downstream_readdatavalid : OUT STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_reset_n : OUT STD_LOGIC;
                    signal nios2_fpu_burst_6_downstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_6_downstream_arbitrator;

component nios2_fpu_burst_6 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_6;

component nios2_fpu_burst_7_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal nios2_fast_fpu_instruction_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fast_fpu_instruction_master_latency_counter : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fpu_burst_7_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_7_upstream_readdatavalid : IN STD_LOGIC;
                    signal nios2_fpu_burst_7_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_nios2_fpu_burst_7_upstream_end_xfer : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register : OUT STD_LOGIC;
                    signal nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream : OUT STD_LOGIC;
                    signal nios2_fpu_burst_7_upstream_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_burst_7_upstream_byteaddress : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal nios2_fpu_burst_7_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_7_upstream_debugaccess : OUT STD_LOGIC;
                    signal nios2_fpu_burst_7_upstream_read : OUT STD_LOGIC;
                    signal nios2_fpu_burst_7_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_7_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_fpu_burst_7_upstream_write : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_7_upstream_arbitrator;

component nios2_fpu_burst_7_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_ipl_memory_s1_end_xfer : IN STD_LOGIC;
                    signal ipl_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_7_downstream_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_burst_7_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_7_downstream_granted_ipl_memory_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_requests_ipl_memory_s1 : IN STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_fpu_burst_7_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_burst_7_downstream_latency_counter : OUT STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_7_downstream_readdatavalid : OUT STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_reset_n : OUT STD_LOGIC;
                    signal nios2_fpu_burst_7_downstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_7_downstream_arbitrator;

component nios2_fpu_burst_7 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_7;

component nios2_fpu_burst_8_upstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (28 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fast_fpu_data_master_debugaccess : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_latency_counter : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_write : IN STD_LOGIC;
                    signal nios2_fast_fpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_8_upstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_8_upstream_readdatavalid : IN STD_LOGIC;
                    signal nios2_fpu_burst_8_upstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_nios2_fpu_burst_8_upstream_end_xfer : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register : OUT STD_LOGIC;
                    signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream : OUT STD_LOGIC;
                    signal nios2_fpu_burst_8_upstream_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_burst_8_upstream_burstcount : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_8_upstream_byteaddress : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal nios2_fpu_burst_8_upstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_8_upstream_debugaccess : OUT STD_LOGIC;
                    signal nios2_fpu_burst_8_upstream_read : OUT STD_LOGIC;
                    signal nios2_fpu_burst_8_upstream_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_8_upstream_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_fpu_burst_8_upstream_write : OUT STD_LOGIC;
                    signal nios2_fpu_burst_8_upstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component nios2_fpu_burst_8_upstream_arbitrator;

component nios2_fpu_burst_8_downstream_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_nios2_fpu_clock_0_in_end_xfer : IN STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_burst_8_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in : IN STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in : IN STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_read_data_valid_nios2_fpu_clock_0_in : IN STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in : IN STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_clock_0_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_clock_0_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_fpu_burst_8_downstream_address_to_slave : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_burst_8_downstream_latency_counter : OUT STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_burst_8_downstream_readdatavalid : OUT STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_reset_n : OUT STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_8_downstream_arbitrator;

component nios2_fpu_burst_8 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal downstream_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal downstream_readdatavalid : IN STD_LOGIC;
                    signal downstream_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal upstream_address : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal upstream_burstcount : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal upstream_debugaccess : IN STD_LOGIC;
                    signal upstream_nativeaddress : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal upstream_read : IN STD_LOGIC;
                    signal upstream_write : IN STD_LOGIC;
                    signal upstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal reg_downstream_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal reg_downstream_arbitrationshare : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_burstcount : OUT STD_LOGIC;
                    signal reg_downstream_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reg_downstream_debugaccess : OUT STD_LOGIC;
                    signal reg_downstream_nativeaddress : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal reg_downstream_read : OUT STD_LOGIC;
                    signal reg_downstream_write : OUT STD_LOGIC;
                    signal reg_downstream_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal upstream_readdatavalid : OUT STD_LOGIC;
                    signal upstream_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_burst_8;

component nios2_fpu_clock_0_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_burst_8_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_8_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_burst_8_downstream_latency_counter : IN STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_nativeaddress : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_burst_8_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_clock_0_in_endofpacket : IN STD_LOGIC;
                    signal nios2_fpu_clock_0_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_clock_0_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_nios2_fpu_clock_0_in_end_xfer : OUT STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in : OUT STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in : OUT STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_read_data_valid_nios2_fpu_clock_0_in : OUT STD_LOGIC;
                    signal nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in : OUT STD_LOGIC;
                    signal nios2_fpu_clock_0_in_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_clock_0_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_clock_0_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal nios2_fpu_clock_0_in_nativeaddress : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal nios2_fpu_clock_0_in_read : OUT STD_LOGIC;
                    signal nios2_fpu_clock_0_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_clock_0_in_reset_n : OUT STD_LOGIC;
                    signal nios2_fpu_clock_0_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal nios2_fpu_clock_0_in_write : OUT STD_LOGIC;
                    signal nios2_fpu_clock_0_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component nios2_fpu_clock_0_in_arbitrator;

component nios2_fpu_clock_0_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_peripheral_bridge_s1_end_xfer : IN STD_LOGIC;
                    signal nios2_fpu_clock_0_out_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_clock_0_out_granted_peripheral_bridge_s1 : IN STD_LOGIC;
                    signal nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1 : IN STD_LOGIC;
                    signal nios2_fpu_clock_0_out_read : IN STD_LOGIC;
                    signal nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1 : IN STD_LOGIC;
                    signal nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1_shift_register : IN STD_LOGIC;
                    signal nios2_fpu_clock_0_out_requests_peripheral_bridge_s1 : IN STD_LOGIC;
                    signal nios2_fpu_clock_0_out_write : IN STD_LOGIC;
                    signal nios2_fpu_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal peripheral_bridge_s1_endofpacket_from_sa : IN STD_LOGIC;
                    signal peripheral_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal peripheral_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal nios2_fpu_clock_0_out_address_to_slave : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_clock_0_out_endofpacket : OUT STD_LOGIC;
                    signal nios2_fpu_clock_0_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal nios2_fpu_clock_0_out_reset_n : OUT STD_LOGIC;
                    signal nios2_fpu_clock_0_out_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_clock_0_out_arbitrator;

component nios2_fpu_clock_0 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component nios2_fpu_clock_0;

component peripheral_bridge_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fpu_clock_0_out_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal nios2_fpu_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal nios2_fpu_clock_0_out_nativeaddress : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal nios2_fpu_clock_0_out_read : IN STD_LOGIC;
                    signal nios2_fpu_clock_0_out_write : IN STD_LOGIC;
                    signal nios2_fpu_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal peripheral_bridge_s1_endofpacket : IN STD_LOGIC;
                    signal peripheral_bridge_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal peripheral_bridge_s1_readdatavalid : IN STD_LOGIC;
                    signal peripheral_bridge_s1_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_peripheral_bridge_s1_end_xfer : OUT STD_LOGIC;
                    signal nios2_fpu_clock_0_out_granted_peripheral_bridge_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1_shift_register : OUT STD_LOGIC;
                    signal nios2_fpu_clock_0_out_requests_peripheral_bridge_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_s1_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal peripheral_bridge_s1_arbiterlock : OUT STD_LOGIC;
                    signal peripheral_bridge_s1_arbiterlock2 : OUT STD_LOGIC;
                    signal peripheral_bridge_s1_burstcount : OUT STD_LOGIC;
                    signal peripheral_bridge_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal peripheral_bridge_s1_chipselect : OUT STD_LOGIC;
                    signal peripheral_bridge_s1_debugaccess : OUT STD_LOGIC;
                    signal peripheral_bridge_s1_endofpacket_from_sa : OUT STD_LOGIC;
                    signal peripheral_bridge_s1_nativeaddress : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal peripheral_bridge_s1_read : OUT STD_LOGIC;
                    signal peripheral_bridge_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal peripheral_bridge_s1_reset_n : OUT STD_LOGIC;
                    signal peripheral_bridge_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal peripheral_bridge_s1_write : OUT STD_LOGIC;
                    signal peripheral_bridge_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component peripheral_bridge_s1_arbitrator;

component peripheral_bridge_m1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_dipsw_s1_end_xfer : IN STD_LOGIC;
                    signal d1_gpio0_s1_end_xfer : IN STD_LOGIC;
                    signal d1_jtag_uart_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                    signal d1_led_s1_end_xfer : IN STD_LOGIC;
                    signal d1_mmcdma_s1_end_xfer : IN STD_LOGIC;
                    signal d1_psw_s1_end_xfer : IN STD_LOGIC;
                    signal d1_spu_s1_end_xfer : IN STD_LOGIC;
                    signal d1_sysid_control_slave_end_xfer : IN STD_LOGIC;
                    signal d1_systimer_s1_end_xfer : IN STD_LOGIC;
                    signal d1_sysuart_s1_end_xfer : IN STD_LOGIC;
                    signal d1_vga_s1_end_xfer : IN STD_LOGIC;
                    signal dipsw_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal gpio0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal led_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal mmcdma_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal mmcdma_s1_wait_counter_eq_0 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                    signal peripheral_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                    signal peripheral_bridge_m1_granted_dipsw_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_granted_gpio0_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal peripheral_bridge_m1_granted_led_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_granted_mmcdma_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_granted_psw_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_granted_spu_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_granted_sysid_control_slave : IN STD_LOGIC;
                    signal peripheral_bridge_m1_granted_systimer_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_granted_sysuart_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_granted_vga_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_dipsw_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_gpio0_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_led_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_mmcdma_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_psw_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_spu_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_sysid_control_slave : IN STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_systimer_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_sysuart_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_vga_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_dipsw_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_gpio0_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_led_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_mmcdma_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_psw_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_spu_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_sysid_control_slave : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_systimer_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_sysuart_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_vga_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_requests_dipsw_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_requests_gpio0_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal peripheral_bridge_m1_requests_led_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_requests_mmcdma_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_requests_psw_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_requests_spu_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_requests_sysid_control_slave : IN STD_LOGIC;
                    signal peripheral_bridge_m1_requests_systimer_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_requests_sysuart_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_requests_vga_s1 : IN STD_LOGIC;
                    signal peripheral_bridge_m1_write : IN STD_LOGIC;
                    signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal psw_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal spu_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal spu_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal sysid_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal systimer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sysuart_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal vga_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal peripheral_bridge_m1_address_to_slave : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal peripheral_bridge_m1_latency_counter : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal peripheral_bridge_m1_readdatavalid : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_waitrequest : OUT STD_LOGIC
                 );
end component peripheral_bridge_m1_arbitrator;

component peripheral_bridge is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal m1_endofpacket : IN STD_LOGIC;
                    signal m1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal m1_readdatavalid : IN STD_LOGIC;
                    signal m1_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal s1_address : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal s1_arbiterlock : IN STD_LOGIC;
                    signal s1_arbiterlock2 : IN STD_LOGIC;
                    signal s1_burstcount : IN STD_LOGIC;
                    signal s1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal s1_chipselect : IN STD_LOGIC;
                    signal s1_debugaccess : IN STD_LOGIC;
                    signal s1_nativeaddress : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal s1_read : IN STD_LOGIC;
                    signal s1_write : IN STD_LOGIC;
                    signal s1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal m1_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal m1_burstcount : OUT STD_LOGIC;
                    signal m1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m1_chipselect : OUT STD_LOGIC;
                    signal m1_debugaccess : OUT STD_LOGIC;
                    signal m1_read : OUT STD_LOGIC;
                    signal m1_write : OUT STD_LOGIC;
                    signal m1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal s1_endofpacket : OUT STD_LOGIC;
                    signal s1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal s1_readdatavalid : OUT STD_LOGIC;
                    signal s1_waitrequest : OUT STD_LOGIC
                 );
end component peripheral_bridge;

component peripheral_bridge_bridge_arbitrator is 
end component peripheral_bridge_bridge_arbitrator;

component psw_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                    signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                    signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read : IN STD_LOGIC;
                    signal peripheral_bridge_m1_write : IN STD_LOGIC;
                    signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal psw_s1_irq : IN STD_LOGIC;
                    signal psw_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_psw_s1_end_xfer : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_granted_psw_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_psw_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_psw_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_requests_psw_s1 : OUT STD_LOGIC;
                    signal psw_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal psw_s1_chipselect : OUT STD_LOGIC;
                    signal psw_s1_irq_from_sa : OUT STD_LOGIC;
                    signal psw_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal psw_s1_reset_n : OUT STD_LOGIC;
                    signal psw_s1_write_n : OUT STD_LOGIC;
                    signal psw_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component psw_s1_arbitrator;

component psw is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal in_port : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component psw;

component sdram_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_0_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal nios2_fpu_burst_0_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fpu_burst_0_downstream_latency_counter : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_1_downstream_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_1_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal nios2_fpu_burst_1_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fpu_burst_1_downstream_latency_counter : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_2_downstream_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_2_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal nios2_fpu_burst_2_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fpu_burst_2_downstream_latency_counter : IN STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_3_downstream_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal nios2_fpu_burst_3_downstream_arbitrationshare : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal nios2_fpu_burst_3_downstream_burstcount : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal nios2_fpu_burst_3_downstream_latency_counter : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_read : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_write : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_s1_readdatavalid : IN STD_LOGIC;
                    signal sdram_s1_waitrequest : IN STD_LOGIC;

                 -- outputs:
                    signal d1_sdram_s1_end_xfer : OUT STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_granted_sdram_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_qualified_request_sdram_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                    signal nios2_fpu_burst_0_downstream_requests_sdram_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_granted_sdram_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_qualified_request_sdram_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                    signal nios2_fpu_burst_1_downstream_requests_sdram_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_granted_sdram_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_qualified_request_sdram_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                    signal nios2_fpu_burst_2_downstream_requests_sdram_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_granted_sdram_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_qualified_request_sdram_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                    signal nios2_fpu_burst_3_downstream_requests_sdram_s1 : OUT STD_LOGIC;
                    signal sdram_s1_address : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal sdram_s1_byteenable_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal sdram_s1_chipselect : OUT STD_LOGIC;
                    signal sdram_s1_read_n : OUT STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_s1_reset_n : OUT STD_LOGIC;
                    signal sdram_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal sdram_s1_write_n : OUT STD_LOGIC;
                    signal sdram_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sdram_s1_arbitrator;

component sdram is 
           port (
                 -- inputs:
                    signal az_addr : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal az_be_n : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal az_cs : IN STD_LOGIC;
                    signal az_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal az_rd_n : IN STD_LOGIC;
                    signal az_wr_n : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal za_data : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal za_valid : OUT STD_LOGIC;
                    signal za_waitrequest : OUT STD_LOGIC;
                    signal zs_addr : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal zs_ba : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_cas_n : OUT STD_LOGIC;
                    signal zs_cke : OUT STD_LOGIC;
                    signal zs_cs_n : OUT STD_LOGIC;
                    signal zs_dq : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal zs_dqm : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_ras_n : OUT STD_LOGIC;
                    signal zs_we_n : OUT STD_LOGIC
                 );
end component sdram;

component spu_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                    signal peripheral_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                    signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read : IN STD_LOGIC;
                    signal peripheral_bridge_m1_write : IN STD_LOGIC;
                    signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal spu_s1_irq : IN STD_LOGIC;
                    signal spu_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal spu_s1_waitrequest : IN STD_LOGIC;

                 -- outputs:
                    signal d1_spu_s1_end_xfer : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_granted_spu_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_spu_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_spu_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_requests_spu_s1 : OUT STD_LOGIC;
                    signal spu_s1_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal spu_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal spu_s1_chipselect : OUT STD_LOGIC;
                    signal spu_s1_irq_from_sa : OUT STD_LOGIC;
                    signal spu_s1_read : OUT STD_LOGIC;
                    signal spu_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal spu_s1_reset : OUT STD_LOGIC;
                    signal spu_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal spu_s1_write : OUT STD_LOGIC;
                    signal spu_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component spu_s1_arbitrator;

component spu_m1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_nios2_fpu_burst_3_upstream_end_xfer : IN STD_LOGIC;
                    signal nios2_fpu_burst_3_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_3_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal spu_m1_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal spu_m1_burstcount : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal spu_m1_granted_nios2_fpu_burst_3_upstream : IN STD_LOGIC;
                    signal spu_m1_qualified_request_nios2_fpu_burst_3_upstream : IN STD_LOGIC;
                    signal spu_m1_read : IN STD_LOGIC;
                    signal spu_m1_read_data_valid_nios2_fpu_burst_3_upstream : IN STD_LOGIC;
                    signal spu_m1_read_data_valid_nios2_fpu_burst_3_upstream_shift_register : IN STD_LOGIC;
                    signal spu_m1_requests_nios2_fpu_burst_3_upstream : IN STD_LOGIC;

                 -- outputs:
                    signal spu_m1_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal spu_m1_latency_counter : OUT STD_LOGIC;
                    signal spu_m1_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal spu_m1_readdatavalid : OUT STD_LOGIC;
                    signal spu_m1_waitrequest : OUT STD_LOGIC
                 );
end component spu_m1_arbitrator;

component spu is 
           port (
                 -- inputs:
                    signal avm_m1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal avm_m1_readdatavalid : IN STD_LOGIC;
                    signal avm_m1_waitrequest : IN STD_LOGIC;
                    signal avs_s1_address : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal avs_s1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal avs_s1_chipselect : IN STD_LOGIC;
                    signal avs_s1_read : IN STD_LOGIC;
                    signal avs_s1_write : IN STD_LOGIC;
                    signal avs_s1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk_128fs : IN STD_LOGIC;
                    signal csi_global_clock : IN STD_LOGIC;
                    signal csi_global_reset : IN STD_LOGIC;
                    signal csi_m1_clock : IN STD_LOGIC;

                 -- outputs:
                    signal AUD_L : OUT STD_LOGIC;
                    signal AUD_R : OUT STD_LOGIC;
                    signal DAC_BCLK : OUT STD_LOGIC;
                    signal DAC_DATA : OUT STD_LOGIC;
                    signal DAC_LRCK : OUT STD_LOGIC;
                    signal SPDIF : OUT STD_LOGIC;
                    signal avm_m1_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal avm_m1_burstcount : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal avm_m1_read : OUT STD_LOGIC;
                    signal avs_s1_irq : OUT STD_LOGIC;
                    signal avs_s1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal avs_s1_waitrequest : OUT STD_LOGIC
                 );
end component spu;

component sysid_control_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                    signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                    signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read : IN STD_LOGIC;
                    signal peripheral_bridge_m1_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sysid_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal d1_sysid_control_slave_end_xfer : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_granted_sysid_control_slave : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_sysid_control_slave : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_sysid_control_slave : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_requests_sysid_control_slave : OUT STD_LOGIC;
                    signal sysid_control_slave_address : OUT STD_LOGIC;
                    signal sysid_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sysid_control_slave_reset_n : OUT STD_LOGIC
                 );
end component sysid_control_slave_arbitrator;

component sysid is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC;
                    signal clock : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sysid;

component systimer_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                    signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                    signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read : IN STD_LOGIC;
                    signal peripheral_bridge_m1_write : IN STD_LOGIC;
                    signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal systimer_s1_irq : IN STD_LOGIC;
                    signal systimer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal d1_systimer_s1_end_xfer : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_granted_systimer_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_systimer_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_systimer_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_requests_systimer_s1 : OUT STD_LOGIC;
                    signal systimer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal systimer_s1_chipselect : OUT STD_LOGIC;
                    signal systimer_s1_irq_from_sa : OUT STD_LOGIC;
                    signal systimer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal systimer_s1_reset_n : OUT STD_LOGIC;
                    signal systimer_s1_write_n : OUT STD_LOGIC;
                    signal systimer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component systimer_s1_arbitrator;

component systimer is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component systimer;

component sysuart_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                    signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                    signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read : IN STD_LOGIC;
                    signal peripheral_bridge_m1_write : IN STD_LOGIC;
                    signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sysuart_s1_dataavailable : IN STD_LOGIC;
                    signal sysuart_s1_irq : IN STD_LOGIC;
                    signal sysuart_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sysuart_s1_readyfordata : IN STD_LOGIC;

                 -- outputs:
                    signal d1_sysuart_s1_end_xfer : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_granted_sysuart_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_sysuart_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_sysuart_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_requests_sysuart_s1 : OUT STD_LOGIC;
                    signal sysuart_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal sysuart_s1_begintransfer : OUT STD_LOGIC;
                    signal sysuart_s1_chipselect : OUT STD_LOGIC;
                    signal sysuart_s1_dataavailable_from_sa : OUT STD_LOGIC;
                    signal sysuart_s1_irq_from_sa : OUT STD_LOGIC;
                    signal sysuart_s1_read_n : OUT STD_LOGIC;
                    signal sysuart_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sysuart_s1_readyfordata_from_sa : OUT STD_LOGIC;
                    signal sysuart_s1_reset_n : OUT STD_LOGIC;
                    signal sysuart_s1_write_n : OUT STD_LOGIC;
                    signal sysuart_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sysuart_s1_arbitrator;

component sysuart is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal begintransfer : IN STD_LOGIC;
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read_n : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal rxd : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal dataavailable : OUT STD_LOGIC;
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readyfordata : OUT STD_LOGIC;
                    signal txd : OUT STD_LOGIC
                 );
end component sysuart;

component vga_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal peripheral_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal peripheral_bridge_m1_burstcount : IN STD_LOGIC;
                    signal peripheral_bridge_m1_chipselect : IN STD_LOGIC;
                    signal peripheral_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal peripheral_bridge_m1_read : IN STD_LOGIC;
                    signal peripheral_bridge_m1_write : IN STD_LOGIC;
                    signal peripheral_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal vga_s1_irq : IN STD_LOGIC;
                    signal vga_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal d1_vga_s1_end_xfer : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_granted_vga_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_qualified_request_vga_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_read_data_valid_vga_s1 : OUT STD_LOGIC;
                    signal peripheral_bridge_m1_requests_vga_s1 : OUT STD_LOGIC;
                    signal vga_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal vga_s1_irq_from_sa : OUT STD_LOGIC;
                    signal vga_s1_read : OUT STD_LOGIC;
                    signal vga_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal vga_s1_write : OUT STD_LOGIC;
                    signal vga_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component vga_s1_arbitrator;

component vga_m1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_nios2_fpu_burst_0_upstream_end_xfer : IN STD_LOGIC;
                    signal nios2_fpu_burst_0_upstream_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal nios2_fpu_burst_0_upstream_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal vga_m1_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal vga_m1_burstcount : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal vga_m1_granted_nios2_fpu_burst_0_upstream : IN STD_LOGIC;
                    signal vga_m1_qualified_request_nios2_fpu_burst_0_upstream : IN STD_LOGIC;
                    signal vga_m1_read : IN STD_LOGIC;
                    signal vga_m1_read_data_valid_nios2_fpu_burst_0_upstream : IN STD_LOGIC;
                    signal vga_m1_read_data_valid_nios2_fpu_burst_0_upstream_shift_register : IN STD_LOGIC;
                    signal vga_m1_requests_nios2_fpu_burst_0_upstream : IN STD_LOGIC;

                 -- outputs:
                    signal vga_m1_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal vga_m1_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal vga_m1_latency_counter : OUT STD_LOGIC;
                    signal vga_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal vga_m1_readdatavalid : OUT STD_LOGIC;
                    signal vga_m1_reset : OUT STD_LOGIC;
                    signal vga_m1_waitrequest : OUT STD_LOGIC
                 );
end component vga_m1_arbitrator;

component vga is 
           port (
                 -- inputs:
                    signal avm_m1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal avm_m1_readdatavalid : IN STD_LOGIC;
                    signal avm_m1_waitrequest : IN STD_LOGIC;
                    signal avs_s1_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal avs_s1_read : IN STD_LOGIC;
                    signal avs_s1_write : IN STD_LOGIC;
                    signal avs_s1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal csi_m1_clk : IN STD_LOGIC;
                    signal csi_m1_reset : IN STD_LOGIC;
                    signal csi_s1_clk : IN STD_LOGIC;
                    signal video_clk : IN STD_LOGIC;

                 -- outputs:
                    signal avm_m1_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal avm_m1_burstcount : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal avm_m1_read : OUT STD_LOGIC;
                    signal avs_s1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal irq_s1 : OUT STD_LOGIC;
                    signal video_bout : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal video_enable : OUT STD_LOGIC;
                    signal video_gout : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal video_hsync_n : OUT STD_LOGIC;
                    signal video_rout : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal video_vsync_n : OUT STD_LOGIC
                 );
end component vga;

component nios2_fpu_reset_peri_clk_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component nios2_fpu_reset_peri_clk_domain_synch_module;

component nios2_fpu_reset_core_clk_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component nios2_fpu_reset_core_clk_domain_synch_module;

                signal core_clk_reset_n :  STD_LOGIC;
                signal d1_dipsw_s1_end_xfer :  STD_LOGIC;
                signal d1_gpio0_s1_end_xfer :  STD_LOGIC;
                signal d1_ipl_memory_s1_end_xfer :  STD_LOGIC;
                signal d1_jtag_uart_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal d1_led_s1_end_xfer :  STD_LOGIC;
                signal d1_mmcdma_s1_end_xfer :  STD_LOGIC;
                signal d1_nios2_fast_fpu_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal d1_nios2_fpu_burst_0_upstream_end_xfer :  STD_LOGIC;
                signal d1_nios2_fpu_burst_1_upstream_end_xfer :  STD_LOGIC;
                signal d1_nios2_fpu_burst_2_upstream_end_xfer :  STD_LOGIC;
                signal d1_nios2_fpu_burst_3_upstream_end_xfer :  STD_LOGIC;
                signal d1_nios2_fpu_burst_4_upstream_end_xfer :  STD_LOGIC;
                signal d1_nios2_fpu_burst_5_upstream_end_xfer :  STD_LOGIC;
                signal d1_nios2_fpu_burst_6_upstream_end_xfer :  STD_LOGIC;
                signal d1_nios2_fpu_burst_7_upstream_end_xfer :  STD_LOGIC;
                signal d1_nios2_fpu_burst_8_upstream_end_xfer :  STD_LOGIC;
                signal d1_nios2_fpu_clock_0_in_end_xfer :  STD_LOGIC;
                signal d1_peripheral_bridge_s1_end_xfer :  STD_LOGIC;
                signal d1_psw_s1_end_xfer :  STD_LOGIC;
                signal d1_sdram_s1_end_xfer :  STD_LOGIC;
                signal d1_spu_s1_end_xfer :  STD_LOGIC;
                signal d1_sysid_control_slave_end_xfer :  STD_LOGIC;
                signal d1_systimer_s1_end_xfer :  STD_LOGIC;
                signal d1_sysuart_s1_end_xfer :  STD_LOGIC;
                signal d1_vga_s1_end_xfer :  STD_LOGIC;
                signal dipsw_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal dipsw_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dipsw_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dipsw_s1_reset_n :  STD_LOGIC;
                signal gpio0_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gpio0_s1_chipselect :  STD_LOGIC;
                signal gpio0_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal gpio0_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal gpio0_s1_reset_n :  STD_LOGIC;
                signal gpio0_s1_write_n :  STD_LOGIC;
                signal gpio0_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_AUD_L_from_the_spu :  STD_LOGIC;
                signal internal_AUD_R_from_the_spu :  STD_LOGIC;
                signal internal_DAC_BCLK_from_the_spu :  STD_LOGIC;
                signal internal_DAC_DATA_from_the_spu :  STD_LOGIC;
                signal internal_DAC_LRCK_from_the_spu :  STD_LOGIC;
                signal internal_MMC_SCK_from_the_mmcdma :  STD_LOGIC;
                signal internal_MMC_SDO_from_the_mmcdma :  STD_LOGIC;
                signal internal_MMC_nCS_from_the_mmcdma :  STD_LOGIC;
                signal internal_SPDIF_from_the_spu :  STD_LOGIC;
                signal internal_out_port_from_the_led :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_txd_from_the_sysuart :  STD_LOGIC;
                signal internal_video_bout_from_the_vga :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal internal_video_enable_from_the_vga :  STD_LOGIC;
                signal internal_video_gout_from_the_vga :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal internal_video_hsync_n_from_the_vga :  STD_LOGIC;
                signal internal_video_rout_from_the_vga :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal internal_video_vsync_n_from_the_vga :  STD_LOGIC;
                signal internal_zs_addr_from_the_sdram :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal internal_zs_ba_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_zs_cas_n_from_the_sdram :  STD_LOGIC;
                signal internal_zs_cke_from_the_sdram :  STD_LOGIC;
                signal internal_zs_cs_n_from_the_sdram :  STD_LOGIC;
                signal internal_zs_dqm_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_zs_ras_n_from_the_sdram :  STD_LOGIC;
                signal internal_zs_we_n_from_the_sdram :  STD_LOGIC;
                signal ipl_memory_s1_address :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal ipl_memory_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ipl_memory_s1_chipselect :  STD_LOGIC;
                signal ipl_memory_s1_clken :  STD_LOGIC;
                signal ipl_memory_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ipl_memory_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ipl_memory_s1_reset :  STD_LOGIC;
                signal ipl_memory_s1_write :  STD_LOGIC;
                signal ipl_memory_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_address :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_chipselect :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_dataavailable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_irq :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_irq_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_read_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_readyfordata :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_reset_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waitrequest :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_write_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal led_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal led_s1_chipselect :  STD_LOGIC;
                signal led_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal led_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal led_s1_reset_n :  STD_LOGIC;
                signal led_s1_write_n :  STD_LOGIC;
                signal led_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal mmcdma_s1_address :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal mmcdma_s1_chipselect :  STD_LOGIC;
                signal mmcdma_s1_irq :  STD_LOGIC;
                signal mmcdma_s1_irq_from_sa :  STD_LOGIC;
                signal mmcdma_s1_read :  STD_LOGIC;
                signal mmcdma_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal mmcdma_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal mmcdma_s1_reset :  STD_LOGIC;
                signal mmcdma_s1_wait_counter_eq_0 :  STD_LOGIC;
                signal mmcdma_s1_write :  STD_LOGIC;
                signal mmcdma_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal module_input69 :  STD_LOGIC;
                signal module_input70 :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_a :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fast_fpu_custom_instruction_master_multi_b :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fast_fpu_custom_instruction_master_multi_c :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fast_fpu_custom_instruction_master_multi_clk :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_clk_en :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_dataa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_custom_instruction_master_multi_datab :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_custom_instruction_master_multi_done :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_estatus :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_ipending :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_custom_instruction_master_multi_n :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal nios2_fast_fpu_custom_instruction_master_multi_readra :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_readrb :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_reset :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_result :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_custom_instruction_master_multi_start :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_status :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_writerc :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_reset_n :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_fpoint_s1 :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0 :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_address :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal nios2_fast_fpu_data_master_address_to_slave :  STD_LOGIC_VECTOR (28 DOWNTO 0);
                signal nios2_fast_fpu_data_master_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fast_fpu_data_master_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_data_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_data_master_dbs_write_16 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fast_fpu_data_master_debugaccess :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_irq :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_data_master_latency_counter :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_read :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_data_master_readdatavalid :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_waitrequest :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_write :  STD_LOGIC;
                signal nios2_fast_fpu_data_master_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_fpoint_s1_clk_en :  STD_LOGIC;
                signal nios2_fast_fpu_fpoint_s1_dataa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_fpoint_s1_datab :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_fpoint_s1_done :  STD_LOGIC;
                signal nios2_fast_fpu_fpoint_s1_done_from_sa :  STD_LOGIC;
                signal nios2_fast_fpu_fpoint_s1_n :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_fpoint_s1_reset :  STD_LOGIC;
                signal nios2_fast_fpu_fpoint_s1_result :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_fpoint_s1_result_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_fpoint_s1_select :  STD_LOGIC;
                signal nios2_fast_fpu_fpoint_s1_start :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_address :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal nios2_fast_fpu_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal nios2_fast_fpu_instruction_master_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fast_fpu_instruction_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_latency_counter :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_read :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_instruction_master_readdatavalid :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream :  STD_LOGIC;
                signal nios2_fast_fpu_instruction_master_waitrequest :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_address :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal nios2_fast_fpu_jtag_debug_module_begintransfer :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fast_fpu_jtag_debug_module_chipselect :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_debugaccess :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_jtag_debug_module_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_jtag_debug_module_resetrequest :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_resetrequest_from_sa :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_write :  STD_LOGIC;
                signal nios2_fast_fpu_jtag_debug_module_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_clk_en :  STD_LOGIC;
                signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_dataa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_datab :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done :  STD_LOGIC;
                signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done_from_sa :  STD_LOGIC;
                signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_n :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_reset :  STD_LOGIC;
                signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select :  STD_LOGIC;
                signal nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_start :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_0_downstream_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_0_downstream_arbitrationshare :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_0_downstream_burstcount :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fpu_burst_0_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_granted_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_latency_counter :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_nativeaddress :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_0_downstream_qualified_request_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1_shift_register :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_0_downstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_requests_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_reset_n :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_byteaddress :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_0_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_1_downstream_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_1_downstream_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_1_downstream_arbitrationshare :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fpu_burst_1_downstream_burstcount :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fpu_burst_1_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_granted_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_latency_counter :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_nativeaddress :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_1_downstream_qualified_request_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1_shift_register :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_1_downstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_requests_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_reset_n :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_1_upstream_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_1_upstream_byteaddress :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal nios2_fpu_burst_1_upstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fpu_burst_1_upstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_1_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_1_upstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_1_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_2_downstream_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_2_downstream_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_2_downstream_arbitrationshare :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fpu_burst_2_downstream_burstcount :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fpu_burst_2_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_granted_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_latency_counter :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_nativeaddress :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_2_downstream_qualified_request_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1_shift_register :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_2_downstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_requests_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_reset_n :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_byteaddress :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_2_upstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_2_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_3_downstream_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_3_downstream_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_3_downstream_arbitrationshare :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_3_downstream_burstcount :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fpu_burst_3_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_granted_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_latency_counter :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_nativeaddress :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_3_downstream_qualified_request_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1_shift_register :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_3_downstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_requests_sdram_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_reset_n :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_byteaddress :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_3_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_4_downstream_address :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_4_downstream_address_to_slave :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_4_downstream_arbitrationshare :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_4_downstream_burstcount :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_4_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_latency_counter :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_nativeaddress :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_4_downstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_reset_n :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_4_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_4_upstream_address :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_4_upstream_byteaddress :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_4_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_4_upstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_4_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_4_upstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_4_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_5_downstream_address :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_5_downstream_address_to_slave :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_5_downstream_arbitrationshare :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_5_downstream_burstcount :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_5_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_latency_counter :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_nativeaddress :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_5_downstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_reset_n :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_5_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_address :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_byteaddress :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_5_upstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_5_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_6_downstream_address :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_6_downstream_address_to_slave :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_6_downstream_arbitrationshare :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_6_downstream_burstcount :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_6_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_latency_counter :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_nativeaddress :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_6_downstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_requests_ipl_memory_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_reset_n :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_address :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_byteaddress :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_6_upstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_6_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_7_downstream_address :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_7_downstream_address_to_slave :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_7_downstream_arbitrationshare :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_7_downstream_burstcount :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_7_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_granted_ipl_memory_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_latency_counter :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_nativeaddress :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_7_downstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_requests_ipl_memory_s1 :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_reset_n :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_7_upstream_address :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_7_upstream_byteaddress :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal nios2_fpu_burst_7_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_7_upstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_7_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_7_upstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_7_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_8_downstream_address :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_8_downstream_address_to_slave :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_8_downstream_arbitrationshare :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_8_downstream_burstcount :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_8_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_latency_counter :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_nativeaddress :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_read_data_valid_nios2_fpu_clock_0_in :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_8_downstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_reset_n :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_8_downstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_address :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_burstcount :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_byteaddress :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_read :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_8_upstream_readdatavalid :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_waitrequest :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_write :  STD_LOGIC;
                signal nios2_fpu_burst_8_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_clock_0_in_address :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_clock_0_in_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_clock_0_in_endofpacket :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_endofpacket_from_sa :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_nativeaddress :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_clock_0_in_read :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_clock_0_in_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_clock_0_in_reset_n :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_waitrequest :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_waitrequest_from_sa :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_write :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_clock_0_out_address :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_clock_0_out_address_to_slave :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_clock_0_out_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal nios2_fpu_clock_0_out_endofpacket :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_granted_peripheral_bridge_s1 :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_nativeaddress :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1 :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_read :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1 :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1_shift_register :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_clock_0_out_requests_peripheral_bridge_s1 :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_reset_n :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_waitrequest :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_write :  STD_LOGIC;
                signal nios2_fpu_clock_0_out_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal peri_clk_reset_n :  STD_LOGIC;
                signal peripheral_bridge_m1_address :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal peripheral_bridge_m1_address_to_slave :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal peripheral_bridge_m1_burstcount :  STD_LOGIC;
                signal peripheral_bridge_m1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal peripheral_bridge_m1_chipselect :  STD_LOGIC;
                signal peripheral_bridge_m1_debugaccess :  STD_LOGIC;
                signal peripheral_bridge_m1_endofpacket :  STD_LOGIC;
                signal peripheral_bridge_m1_granted_dipsw_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_granted_gpio0_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal peripheral_bridge_m1_granted_led_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_granted_mmcdma_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_granted_psw_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_granted_spu_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_granted_sysid_control_slave :  STD_LOGIC;
                signal peripheral_bridge_m1_granted_systimer_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_granted_sysuart_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_granted_vga_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_latency_counter :  STD_LOGIC;
                signal peripheral_bridge_m1_qualified_request_dipsw_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_qualified_request_gpio0_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal peripheral_bridge_m1_qualified_request_led_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_qualified_request_mmcdma_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_qualified_request_psw_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_qualified_request_spu_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_qualified_request_sysid_control_slave :  STD_LOGIC;
                signal peripheral_bridge_m1_qualified_request_systimer_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_qualified_request_sysuart_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_qualified_request_vga_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_read :  STD_LOGIC;
                signal peripheral_bridge_m1_read_data_valid_dipsw_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_read_data_valid_gpio0_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal peripheral_bridge_m1_read_data_valid_led_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_read_data_valid_mmcdma_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_read_data_valid_psw_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_read_data_valid_spu_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_read_data_valid_sysid_control_slave :  STD_LOGIC;
                signal peripheral_bridge_m1_read_data_valid_systimer_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_read_data_valid_sysuart_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_read_data_valid_vga_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal peripheral_bridge_m1_readdatavalid :  STD_LOGIC;
                signal peripheral_bridge_m1_requests_dipsw_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_requests_gpio0_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal peripheral_bridge_m1_requests_led_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_requests_mmcdma_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_requests_psw_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_requests_spu_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_requests_sysid_control_slave :  STD_LOGIC;
                signal peripheral_bridge_m1_requests_systimer_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_requests_sysuart_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_requests_vga_s1 :  STD_LOGIC;
                signal peripheral_bridge_m1_waitrequest :  STD_LOGIC;
                signal peripheral_bridge_m1_write :  STD_LOGIC;
                signal peripheral_bridge_m1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal peripheral_bridge_s1_address :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal peripheral_bridge_s1_arbiterlock :  STD_LOGIC;
                signal peripheral_bridge_s1_arbiterlock2 :  STD_LOGIC;
                signal peripheral_bridge_s1_burstcount :  STD_LOGIC;
                signal peripheral_bridge_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal peripheral_bridge_s1_chipselect :  STD_LOGIC;
                signal peripheral_bridge_s1_debugaccess :  STD_LOGIC;
                signal peripheral_bridge_s1_endofpacket :  STD_LOGIC;
                signal peripheral_bridge_s1_endofpacket_from_sa :  STD_LOGIC;
                signal peripheral_bridge_s1_nativeaddress :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal peripheral_bridge_s1_read :  STD_LOGIC;
                signal peripheral_bridge_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal peripheral_bridge_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal peripheral_bridge_s1_readdatavalid :  STD_LOGIC;
                signal peripheral_bridge_s1_reset_n :  STD_LOGIC;
                signal peripheral_bridge_s1_waitrequest :  STD_LOGIC;
                signal peripheral_bridge_s1_waitrequest_from_sa :  STD_LOGIC;
                signal peripheral_bridge_s1_write :  STD_LOGIC;
                signal peripheral_bridge_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal psw_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal psw_s1_chipselect :  STD_LOGIC;
                signal psw_s1_irq :  STD_LOGIC;
                signal psw_s1_irq_from_sa :  STD_LOGIC;
                signal psw_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal psw_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal psw_s1_reset_n :  STD_LOGIC;
                signal psw_s1_write_n :  STD_LOGIC;
                signal psw_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal reset_n_sources :  STD_LOGIC;
                signal sdram_s1_address :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal sdram_s1_byteenable_n :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_s1_chipselect :  STD_LOGIC;
                signal sdram_s1_read_n :  STD_LOGIC;
                signal sdram_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sdram_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sdram_s1_readdatavalid :  STD_LOGIC;
                signal sdram_s1_reset_n :  STD_LOGIC;
                signal sdram_s1_waitrequest :  STD_LOGIC;
                signal sdram_s1_waitrequest_from_sa :  STD_LOGIC;
                signal sdram_s1_write_n :  STD_LOGIC;
                signal sdram_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal spu_m1_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal spu_m1_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal spu_m1_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal spu_m1_granted_nios2_fpu_burst_3_upstream :  STD_LOGIC;
                signal spu_m1_latency_counter :  STD_LOGIC;
                signal spu_m1_qualified_request_nios2_fpu_burst_3_upstream :  STD_LOGIC;
                signal spu_m1_read :  STD_LOGIC;
                signal spu_m1_read_data_valid_nios2_fpu_burst_3_upstream :  STD_LOGIC;
                signal spu_m1_read_data_valid_nios2_fpu_burst_3_upstream_shift_register :  STD_LOGIC;
                signal spu_m1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal spu_m1_readdatavalid :  STD_LOGIC;
                signal spu_m1_requests_nios2_fpu_burst_3_upstream :  STD_LOGIC;
                signal spu_m1_waitrequest :  STD_LOGIC;
                signal spu_s1_address :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal spu_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal spu_s1_chipselect :  STD_LOGIC;
                signal spu_s1_irq :  STD_LOGIC;
                signal spu_s1_irq_from_sa :  STD_LOGIC;
                signal spu_s1_read :  STD_LOGIC;
                signal spu_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal spu_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal spu_s1_reset :  STD_LOGIC;
                signal spu_s1_waitrequest :  STD_LOGIC;
                signal spu_s1_waitrequest_from_sa :  STD_LOGIC;
                signal spu_s1_write :  STD_LOGIC;
                signal spu_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sysid_control_slave_address :  STD_LOGIC;
                signal sysid_control_slave_clock :  STD_LOGIC;
                signal sysid_control_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sysid_control_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sysid_control_slave_reset_n :  STD_LOGIC;
                signal systimer_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal systimer_s1_chipselect :  STD_LOGIC;
                signal systimer_s1_irq :  STD_LOGIC;
                signal systimer_s1_irq_from_sa :  STD_LOGIC;
                signal systimer_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal systimer_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal systimer_s1_reset_n :  STD_LOGIC;
                signal systimer_s1_write_n :  STD_LOGIC;
                signal systimer_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sysuart_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sysuart_s1_begintransfer :  STD_LOGIC;
                signal sysuart_s1_chipselect :  STD_LOGIC;
                signal sysuart_s1_dataavailable :  STD_LOGIC;
                signal sysuart_s1_dataavailable_from_sa :  STD_LOGIC;
                signal sysuart_s1_irq :  STD_LOGIC;
                signal sysuart_s1_irq_from_sa :  STD_LOGIC;
                signal sysuart_s1_read_n :  STD_LOGIC;
                signal sysuart_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sysuart_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sysuart_s1_readyfordata :  STD_LOGIC;
                signal sysuart_s1_readyfordata_from_sa :  STD_LOGIC;
                signal sysuart_s1_reset_n :  STD_LOGIC;
                signal sysuart_s1_write_n :  STD_LOGIC;
                signal sysuart_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal vga_m1_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal vga_m1_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal vga_m1_burstcount :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal vga_m1_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal vga_m1_granted_nios2_fpu_burst_0_upstream :  STD_LOGIC;
                signal vga_m1_latency_counter :  STD_LOGIC;
                signal vga_m1_qualified_request_nios2_fpu_burst_0_upstream :  STD_LOGIC;
                signal vga_m1_read :  STD_LOGIC;
                signal vga_m1_read_data_valid_nios2_fpu_burst_0_upstream :  STD_LOGIC;
                signal vga_m1_read_data_valid_nios2_fpu_burst_0_upstream_shift_register :  STD_LOGIC;
                signal vga_m1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal vga_m1_readdatavalid :  STD_LOGIC;
                signal vga_m1_requests_nios2_fpu_burst_0_upstream :  STD_LOGIC;
                signal vga_m1_reset :  STD_LOGIC;
                signal vga_m1_waitrequest :  STD_LOGIC;
                signal vga_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal vga_s1_irq :  STD_LOGIC;
                signal vga_s1_irq_from_sa :  STD_LOGIC;
                signal vga_s1_read :  STD_LOGIC;
                signal vga_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal vga_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal vga_s1_write :  STD_LOGIC;
                signal vga_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);

begin

  --the_dipsw_s1, which is an e_instance
  the_dipsw_s1 : dipsw_s1_arbitrator
    port map(
      d1_dipsw_s1_end_xfer => d1_dipsw_s1_end_xfer,
      dipsw_s1_address => dipsw_s1_address,
      dipsw_s1_readdata_from_sa => dipsw_s1_readdata_from_sa,
      dipsw_s1_reset_n => dipsw_s1_reset_n,
      peripheral_bridge_m1_granted_dipsw_s1 => peripheral_bridge_m1_granted_dipsw_s1,
      peripheral_bridge_m1_qualified_request_dipsw_s1 => peripheral_bridge_m1_qualified_request_dipsw_s1,
      peripheral_bridge_m1_read_data_valid_dipsw_s1 => peripheral_bridge_m1_read_data_valid_dipsw_s1,
      peripheral_bridge_m1_requests_dipsw_s1 => peripheral_bridge_m1_requests_dipsw_s1,
      clk => peri_clk,
      dipsw_s1_readdata => dipsw_s1_readdata,
      peripheral_bridge_m1_address_to_slave => peripheral_bridge_m1_address_to_slave,
      peripheral_bridge_m1_burstcount => peripheral_bridge_m1_burstcount,
      peripheral_bridge_m1_chipselect => peripheral_bridge_m1_chipselect,
      peripheral_bridge_m1_latency_counter => peripheral_bridge_m1_latency_counter,
      peripheral_bridge_m1_read => peripheral_bridge_m1_read,
      peripheral_bridge_m1_write => peripheral_bridge_m1_write,
      reset_n => peri_clk_reset_n
    );


  --the_dipsw, which is an e_ptf_instance
  the_dipsw : dipsw
    port map(
      readdata => dipsw_s1_readdata,
      address => dipsw_s1_address,
      clk => peri_clk,
      in_port => in_port_to_the_dipsw,
      reset_n => dipsw_s1_reset_n
    );


  --the_gpio0_s1, which is an e_instance
  the_gpio0_s1 : gpio0_s1_arbitrator
    port map(
      d1_gpio0_s1_end_xfer => d1_gpio0_s1_end_xfer,
      gpio0_s1_address => gpio0_s1_address,
      gpio0_s1_chipselect => gpio0_s1_chipselect,
      gpio0_s1_readdata_from_sa => gpio0_s1_readdata_from_sa,
      gpio0_s1_reset_n => gpio0_s1_reset_n,
      gpio0_s1_write_n => gpio0_s1_write_n,
      gpio0_s1_writedata => gpio0_s1_writedata,
      peripheral_bridge_m1_granted_gpio0_s1 => peripheral_bridge_m1_granted_gpio0_s1,
      peripheral_bridge_m1_qualified_request_gpio0_s1 => peripheral_bridge_m1_qualified_request_gpio0_s1,
      peripheral_bridge_m1_read_data_valid_gpio0_s1 => peripheral_bridge_m1_read_data_valid_gpio0_s1,
      peripheral_bridge_m1_requests_gpio0_s1 => peripheral_bridge_m1_requests_gpio0_s1,
      clk => peri_clk,
      gpio0_s1_readdata => gpio0_s1_readdata,
      peripheral_bridge_m1_address_to_slave => peripheral_bridge_m1_address_to_slave,
      peripheral_bridge_m1_burstcount => peripheral_bridge_m1_burstcount,
      peripheral_bridge_m1_chipselect => peripheral_bridge_m1_chipselect,
      peripheral_bridge_m1_latency_counter => peripheral_bridge_m1_latency_counter,
      peripheral_bridge_m1_read => peripheral_bridge_m1_read,
      peripheral_bridge_m1_write => peripheral_bridge_m1_write,
      peripheral_bridge_m1_writedata => peripheral_bridge_m1_writedata,
      reset_n => peri_clk_reset_n
    );


  --the_gpio0, which is an e_ptf_instance
  the_gpio0 : gpio0
    port map(
      bidir_port => bidir_port_to_and_from_the_gpio0,
      readdata => gpio0_s1_readdata,
      address => gpio0_s1_address,
      chipselect => gpio0_s1_chipselect,
      clk => peri_clk,
      reset_n => gpio0_s1_reset_n,
      write_n => gpio0_s1_write_n,
      writedata => gpio0_s1_writedata
    );


  --the_ipl_memory_s1, which is an e_instance
  the_ipl_memory_s1 : ipl_memory_s1_arbitrator
    port map(
      d1_ipl_memory_s1_end_xfer => d1_ipl_memory_s1_end_xfer,
      ipl_memory_s1_address => ipl_memory_s1_address,
      ipl_memory_s1_byteenable => ipl_memory_s1_byteenable,
      ipl_memory_s1_chipselect => ipl_memory_s1_chipselect,
      ipl_memory_s1_clken => ipl_memory_s1_clken,
      ipl_memory_s1_readdata_from_sa => ipl_memory_s1_readdata_from_sa,
      ipl_memory_s1_reset => ipl_memory_s1_reset,
      ipl_memory_s1_write => ipl_memory_s1_write,
      ipl_memory_s1_writedata => ipl_memory_s1_writedata,
      nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 => nios2_fpu_burst_6_downstream_granted_ipl_memory_s1,
      nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1 => nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1,
      nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1 => nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1,
      nios2_fpu_burst_6_downstream_requests_ipl_memory_s1 => nios2_fpu_burst_6_downstream_requests_ipl_memory_s1,
      nios2_fpu_burst_7_downstream_granted_ipl_memory_s1 => nios2_fpu_burst_7_downstream_granted_ipl_memory_s1,
      nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1 => nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1,
      nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1 => nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1,
      nios2_fpu_burst_7_downstream_requests_ipl_memory_s1 => nios2_fpu_burst_7_downstream_requests_ipl_memory_s1,
      clk => core_clk,
      ipl_memory_s1_readdata => ipl_memory_s1_readdata,
      nios2_fpu_burst_6_downstream_address_to_slave => nios2_fpu_burst_6_downstream_address_to_slave,
      nios2_fpu_burst_6_downstream_arbitrationshare => nios2_fpu_burst_6_downstream_arbitrationshare,
      nios2_fpu_burst_6_downstream_burstcount => nios2_fpu_burst_6_downstream_burstcount,
      nios2_fpu_burst_6_downstream_byteenable => nios2_fpu_burst_6_downstream_byteenable,
      nios2_fpu_burst_6_downstream_latency_counter => nios2_fpu_burst_6_downstream_latency_counter,
      nios2_fpu_burst_6_downstream_read => nios2_fpu_burst_6_downstream_read,
      nios2_fpu_burst_6_downstream_write => nios2_fpu_burst_6_downstream_write,
      nios2_fpu_burst_6_downstream_writedata => nios2_fpu_burst_6_downstream_writedata,
      nios2_fpu_burst_7_downstream_address_to_slave => nios2_fpu_burst_7_downstream_address_to_slave,
      nios2_fpu_burst_7_downstream_arbitrationshare => nios2_fpu_burst_7_downstream_arbitrationshare,
      nios2_fpu_burst_7_downstream_burstcount => nios2_fpu_burst_7_downstream_burstcount,
      nios2_fpu_burst_7_downstream_byteenable => nios2_fpu_burst_7_downstream_byteenable,
      nios2_fpu_burst_7_downstream_latency_counter => nios2_fpu_burst_7_downstream_latency_counter,
      nios2_fpu_burst_7_downstream_read => nios2_fpu_burst_7_downstream_read,
      nios2_fpu_burst_7_downstream_write => nios2_fpu_burst_7_downstream_write,
      nios2_fpu_burst_7_downstream_writedata => nios2_fpu_burst_7_downstream_writedata,
      reset_n => core_clk_reset_n
    );


  --the_ipl_memory, which is an e_ptf_instance
  the_ipl_memory : ipl_memory
    port map(
      readdata => ipl_memory_s1_readdata,
      address => ipl_memory_s1_address,
      byteenable => ipl_memory_s1_byteenable,
      chipselect => ipl_memory_s1_chipselect,
      clk => core_clk,
      clken => ipl_memory_s1_clken,
      reset => ipl_memory_s1_reset,
      write => ipl_memory_s1_write,
      writedata => ipl_memory_s1_writedata
    );


  --the_jtag_uart_avalon_jtag_slave, which is an e_instance
  the_jtag_uart_avalon_jtag_slave : jtag_uart_avalon_jtag_slave_arbitrator
    port map(
      d1_jtag_uart_avalon_jtag_slave_end_xfer => d1_jtag_uart_avalon_jtag_slave_end_xfer,
      jtag_uart_avalon_jtag_slave_address => jtag_uart_avalon_jtag_slave_address,
      jtag_uart_avalon_jtag_slave_chipselect => jtag_uart_avalon_jtag_slave_chipselect,
      jtag_uart_avalon_jtag_slave_dataavailable_from_sa => jtag_uart_avalon_jtag_slave_dataavailable_from_sa,
      jtag_uart_avalon_jtag_slave_irq_from_sa => jtag_uart_avalon_jtag_slave_irq_from_sa,
      jtag_uart_avalon_jtag_slave_read_n => jtag_uart_avalon_jtag_slave_read_n,
      jtag_uart_avalon_jtag_slave_readdata_from_sa => jtag_uart_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_avalon_jtag_slave_readyfordata_from_sa => jtag_uart_avalon_jtag_slave_readyfordata_from_sa,
      jtag_uart_avalon_jtag_slave_reset_n => jtag_uart_avalon_jtag_slave_reset_n,
      jtag_uart_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
      jtag_uart_avalon_jtag_slave_write_n => jtag_uart_avalon_jtag_slave_write_n,
      jtag_uart_avalon_jtag_slave_writedata => jtag_uart_avalon_jtag_slave_writedata,
      peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave => peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave,
      peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave => peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave,
      peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave => peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave,
      peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave => peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave,
      clk => peri_clk,
      jtag_uart_avalon_jtag_slave_dataavailable => jtag_uart_avalon_jtag_slave_dataavailable,
      jtag_uart_avalon_jtag_slave_irq => jtag_uart_avalon_jtag_slave_irq,
      jtag_uart_avalon_jtag_slave_readdata => jtag_uart_avalon_jtag_slave_readdata,
      jtag_uart_avalon_jtag_slave_readyfordata => jtag_uart_avalon_jtag_slave_readyfordata,
      jtag_uart_avalon_jtag_slave_waitrequest => jtag_uart_avalon_jtag_slave_waitrequest,
      peripheral_bridge_m1_address_to_slave => peripheral_bridge_m1_address_to_slave,
      peripheral_bridge_m1_burstcount => peripheral_bridge_m1_burstcount,
      peripheral_bridge_m1_chipselect => peripheral_bridge_m1_chipselect,
      peripheral_bridge_m1_latency_counter => peripheral_bridge_m1_latency_counter,
      peripheral_bridge_m1_read => peripheral_bridge_m1_read,
      peripheral_bridge_m1_write => peripheral_bridge_m1_write,
      peripheral_bridge_m1_writedata => peripheral_bridge_m1_writedata,
      reset_n => peri_clk_reset_n
    );


  --the_jtag_uart, which is an e_ptf_instance
  the_jtag_uart : jtag_uart
    port map(
      av_irq => jtag_uart_avalon_jtag_slave_irq,
      av_readdata => jtag_uart_avalon_jtag_slave_readdata,
      av_waitrequest => jtag_uart_avalon_jtag_slave_waitrequest,
      dataavailable => jtag_uart_avalon_jtag_slave_dataavailable,
      readyfordata => jtag_uart_avalon_jtag_slave_readyfordata,
      av_address => jtag_uart_avalon_jtag_slave_address,
      av_chipselect => jtag_uart_avalon_jtag_slave_chipselect,
      av_read_n => jtag_uart_avalon_jtag_slave_read_n,
      av_write_n => jtag_uart_avalon_jtag_slave_write_n,
      av_writedata => jtag_uart_avalon_jtag_slave_writedata,
      clk => peri_clk,
      rst_n => jtag_uart_avalon_jtag_slave_reset_n
    );


  --the_led_s1, which is an e_instance
  the_led_s1 : led_s1_arbitrator
    port map(
      d1_led_s1_end_xfer => d1_led_s1_end_xfer,
      led_s1_address => led_s1_address,
      led_s1_chipselect => led_s1_chipselect,
      led_s1_readdata_from_sa => led_s1_readdata_from_sa,
      led_s1_reset_n => led_s1_reset_n,
      led_s1_write_n => led_s1_write_n,
      led_s1_writedata => led_s1_writedata,
      peripheral_bridge_m1_granted_led_s1 => peripheral_bridge_m1_granted_led_s1,
      peripheral_bridge_m1_qualified_request_led_s1 => peripheral_bridge_m1_qualified_request_led_s1,
      peripheral_bridge_m1_read_data_valid_led_s1 => peripheral_bridge_m1_read_data_valid_led_s1,
      peripheral_bridge_m1_requests_led_s1 => peripheral_bridge_m1_requests_led_s1,
      clk => peri_clk,
      led_s1_readdata => led_s1_readdata,
      peripheral_bridge_m1_address_to_slave => peripheral_bridge_m1_address_to_slave,
      peripheral_bridge_m1_burstcount => peripheral_bridge_m1_burstcount,
      peripheral_bridge_m1_chipselect => peripheral_bridge_m1_chipselect,
      peripheral_bridge_m1_latency_counter => peripheral_bridge_m1_latency_counter,
      peripheral_bridge_m1_read => peripheral_bridge_m1_read,
      peripheral_bridge_m1_write => peripheral_bridge_m1_write,
      peripheral_bridge_m1_writedata => peripheral_bridge_m1_writedata,
      reset_n => peri_clk_reset_n
    );


  --the_led, which is an e_ptf_instance
  the_led : led
    port map(
      out_port => internal_out_port_from_the_led,
      readdata => led_s1_readdata,
      address => led_s1_address,
      chipselect => led_s1_chipselect,
      clk => peri_clk,
      reset_n => led_s1_reset_n,
      write_n => led_s1_write_n,
      writedata => led_s1_writedata
    );


  --the_mmcdma_s1, which is an e_instance
  the_mmcdma_s1 : mmcdma_s1_arbitrator
    port map(
      d1_mmcdma_s1_end_xfer => d1_mmcdma_s1_end_xfer,
      mmcdma_s1_address => mmcdma_s1_address,
      mmcdma_s1_chipselect => mmcdma_s1_chipselect,
      mmcdma_s1_irq_from_sa => mmcdma_s1_irq_from_sa,
      mmcdma_s1_read => mmcdma_s1_read,
      mmcdma_s1_readdata_from_sa => mmcdma_s1_readdata_from_sa,
      mmcdma_s1_reset => mmcdma_s1_reset,
      mmcdma_s1_wait_counter_eq_0 => mmcdma_s1_wait_counter_eq_0,
      mmcdma_s1_write => mmcdma_s1_write,
      mmcdma_s1_writedata => mmcdma_s1_writedata,
      peripheral_bridge_m1_granted_mmcdma_s1 => peripheral_bridge_m1_granted_mmcdma_s1,
      peripheral_bridge_m1_qualified_request_mmcdma_s1 => peripheral_bridge_m1_qualified_request_mmcdma_s1,
      peripheral_bridge_m1_read_data_valid_mmcdma_s1 => peripheral_bridge_m1_read_data_valid_mmcdma_s1,
      peripheral_bridge_m1_requests_mmcdma_s1 => peripheral_bridge_m1_requests_mmcdma_s1,
      clk => peri_clk,
      mmcdma_s1_irq => mmcdma_s1_irq,
      mmcdma_s1_readdata => mmcdma_s1_readdata,
      peripheral_bridge_m1_address_to_slave => peripheral_bridge_m1_address_to_slave,
      peripheral_bridge_m1_burstcount => peripheral_bridge_m1_burstcount,
      peripheral_bridge_m1_chipselect => peripheral_bridge_m1_chipselect,
      peripheral_bridge_m1_latency_counter => peripheral_bridge_m1_latency_counter,
      peripheral_bridge_m1_read => peripheral_bridge_m1_read,
      peripheral_bridge_m1_write => peripheral_bridge_m1_write,
      peripheral_bridge_m1_writedata => peripheral_bridge_m1_writedata,
      reset_n => peri_clk_reset_n
    );


  --the_mmcdma, which is an e_ptf_instance
  the_mmcdma : mmcdma
    port map(
      MMC_SCK => internal_MMC_SCK_from_the_mmcdma,
      MMC_SDO => internal_MMC_SDO_from_the_mmcdma,
      MMC_nCS => internal_MMC_nCS_from_the_mmcdma,
      irq => mmcdma_s1_irq,
      readdata => mmcdma_s1_readdata,
      MMC_CD => MMC_CD_to_the_mmcdma,
      MMC_SDI => MMC_SDI_to_the_mmcdma,
      MMC_WP => MMC_WP_to_the_mmcdma,
      address => mmcdma_s1_address,
      chipselect => mmcdma_s1_chipselect,
      clk => peri_clk,
      read => mmcdma_s1_read,
      reset => mmcdma_s1_reset,
      write => mmcdma_s1_write,
      writedata => mmcdma_s1_writedata
    );


  --the_nios2_fast_fpu_jtag_debug_module, which is an e_instance
  the_nios2_fast_fpu_jtag_debug_module : nios2_fast_fpu_jtag_debug_module_arbitrator
    port map(
      d1_nios2_fast_fpu_jtag_debug_module_end_xfer => d1_nios2_fast_fpu_jtag_debug_module_end_xfer,
      nios2_fast_fpu_jtag_debug_module_address => nios2_fast_fpu_jtag_debug_module_address,
      nios2_fast_fpu_jtag_debug_module_begintransfer => nios2_fast_fpu_jtag_debug_module_begintransfer,
      nios2_fast_fpu_jtag_debug_module_byteenable => nios2_fast_fpu_jtag_debug_module_byteenable,
      nios2_fast_fpu_jtag_debug_module_chipselect => nios2_fast_fpu_jtag_debug_module_chipselect,
      nios2_fast_fpu_jtag_debug_module_debugaccess => nios2_fast_fpu_jtag_debug_module_debugaccess,
      nios2_fast_fpu_jtag_debug_module_readdata_from_sa => nios2_fast_fpu_jtag_debug_module_readdata_from_sa,
      nios2_fast_fpu_jtag_debug_module_resetrequest_from_sa => nios2_fast_fpu_jtag_debug_module_resetrequest_from_sa,
      nios2_fast_fpu_jtag_debug_module_write => nios2_fast_fpu_jtag_debug_module_write,
      nios2_fast_fpu_jtag_debug_module_writedata => nios2_fast_fpu_jtag_debug_module_writedata,
      nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module,
      nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module,
      nios2_fpu_burst_4_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_4_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module,
      nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module,
      nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module,
      nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module,
      nios2_fpu_burst_5_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_5_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module,
      nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module,
      clk => core_clk,
      nios2_fast_fpu_jtag_debug_module_readdata => nios2_fast_fpu_jtag_debug_module_readdata,
      nios2_fast_fpu_jtag_debug_module_resetrequest => nios2_fast_fpu_jtag_debug_module_resetrequest,
      nios2_fpu_burst_4_downstream_address_to_slave => nios2_fpu_burst_4_downstream_address_to_slave,
      nios2_fpu_burst_4_downstream_arbitrationshare => nios2_fpu_burst_4_downstream_arbitrationshare,
      nios2_fpu_burst_4_downstream_burstcount => nios2_fpu_burst_4_downstream_burstcount,
      nios2_fpu_burst_4_downstream_byteenable => nios2_fpu_burst_4_downstream_byteenable,
      nios2_fpu_burst_4_downstream_debugaccess => nios2_fpu_burst_4_downstream_debugaccess,
      nios2_fpu_burst_4_downstream_latency_counter => nios2_fpu_burst_4_downstream_latency_counter,
      nios2_fpu_burst_4_downstream_read => nios2_fpu_burst_4_downstream_read,
      nios2_fpu_burst_4_downstream_write => nios2_fpu_burst_4_downstream_write,
      nios2_fpu_burst_4_downstream_writedata => nios2_fpu_burst_4_downstream_writedata,
      nios2_fpu_burst_5_downstream_address_to_slave => nios2_fpu_burst_5_downstream_address_to_slave,
      nios2_fpu_burst_5_downstream_arbitrationshare => nios2_fpu_burst_5_downstream_arbitrationshare,
      nios2_fpu_burst_5_downstream_burstcount => nios2_fpu_burst_5_downstream_burstcount,
      nios2_fpu_burst_5_downstream_byteenable => nios2_fpu_burst_5_downstream_byteenable,
      nios2_fpu_burst_5_downstream_debugaccess => nios2_fpu_burst_5_downstream_debugaccess,
      nios2_fpu_burst_5_downstream_latency_counter => nios2_fpu_burst_5_downstream_latency_counter,
      nios2_fpu_burst_5_downstream_read => nios2_fpu_burst_5_downstream_read,
      nios2_fpu_burst_5_downstream_write => nios2_fpu_burst_5_downstream_write,
      nios2_fpu_burst_5_downstream_writedata => nios2_fpu_burst_5_downstream_writedata,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fast_fpu_custom_instruction_master, which is an e_instance
  the_nios2_fast_fpu_custom_instruction_master : nios2_fast_fpu_custom_instruction_master_arbitrator
    port map(
      nios2_fast_fpu_custom_instruction_master_multi_done => nios2_fast_fpu_custom_instruction_master_multi_done,
      nios2_fast_fpu_custom_instruction_master_multi_result => nios2_fast_fpu_custom_instruction_master_multi_result,
      nios2_fast_fpu_custom_instruction_master_reset_n => nios2_fast_fpu_custom_instruction_master_reset_n,
      nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_fpoint_s1 => nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_fpoint_s1,
      nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0 => nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0,
      nios2_fast_fpu_fpoint_s1_select => nios2_fast_fpu_fpoint_s1_select,
      nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select,
      clk => core_clk,
      nios2_fast_fpu_custom_instruction_master_multi_n => nios2_fast_fpu_custom_instruction_master_multi_n,
      nios2_fast_fpu_custom_instruction_master_multi_start => nios2_fast_fpu_custom_instruction_master_multi_start,
      nios2_fast_fpu_fpoint_s1_done_from_sa => nios2_fast_fpu_fpoint_s1_done_from_sa,
      nios2_fast_fpu_fpoint_s1_result_from_sa => nios2_fast_fpu_fpoint_s1_result_from_sa,
      nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done_from_sa => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done_from_sa,
      nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result_from_sa => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result_from_sa,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fast_fpu_data_master, which is an e_instance
  the_nios2_fast_fpu_data_master : nios2_fast_fpu_data_master_arbitrator
    port map(
      nios2_fast_fpu_data_master_address_to_slave => nios2_fast_fpu_data_master_address_to_slave,
      nios2_fast_fpu_data_master_dbs_address => nios2_fast_fpu_data_master_dbs_address,
      nios2_fast_fpu_data_master_dbs_write_16 => nios2_fast_fpu_data_master_dbs_write_16,
      nios2_fast_fpu_data_master_irq => nios2_fast_fpu_data_master_irq,
      nios2_fast_fpu_data_master_latency_counter => nios2_fast_fpu_data_master_latency_counter,
      nios2_fast_fpu_data_master_readdata => nios2_fast_fpu_data_master_readdata,
      nios2_fast_fpu_data_master_readdatavalid => nios2_fast_fpu_data_master_readdatavalid,
      nios2_fast_fpu_data_master_waitrequest => nios2_fast_fpu_data_master_waitrequest,
      clk => core_clk,
      core_clk => core_clk,
      core_clk_reset_n => core_clk_reset_n,
      d1_nios2_fpu_burst_2_upstream_end_xfer => d1_nios2_fpu_burst_2_upstream_end_xfer,
      d1_nios2_fpu_burst_5_upstream_end_xfer => d1_nios2_fpu_burst_5_upstream_end_xfer,
      d1_nios2_fpu_burst_6_upstream_end_xfer => d1_nios2_fpu_burst_6_upstream_end_xfer,
      d1_nios2_fpu_burst_8_upstream_end_xfer => d1_nios2_fpu_burst_8_upstream_end_xfer,
      jtag_uart_avalon_jtag_slave_irq_from_sa => jtag_uart_avalon_jtag_slave_irq_from_sa,
      mmcdma_s1_irq_from_sa => mmcdma_s1_irq_from_sa,
      nios2_fast_fpu_data_master_address => nios2_fast_fpu_data_master_address,
      nios2_fast_fpu_data_master_burstcount => nios2_fast_fpu_data_master_burstcount,
      nios2_fast_fpu_data_master_byteenable => nios2_fast_fpu_data_master_byteenable,
      nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream => nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream,
      nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream => nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream,
      nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream => nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream,
      nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream => nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream,
      nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream => nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream,
      nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream => nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream,
      nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream => nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream,
      nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream => nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream,
      nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream => nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream,
      nios2_fast_fpu_data_master_read => nios2_fast_fpu_data_master_read,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register,
      nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream => nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream,
      nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream => nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream,
      nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream => nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream,
      nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream => nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream,
      nios2_fast_fpu_data_master_write => nios2_fast_fpu_data_master_write,
      nios2_fast_fpu_data_master_writedata => nios2_fast_fpu_data_master_writedata,
      nios2_fpu_burst_2_upstream_readdata_from_sa => nios2_fpu_burst_2_upstream_readdata_from_sa,
      nios2_fpu_burst_2_upstream_waitrequest_from_sa => nios2_fpu_burst_2_upstream_waitrequest_from_sa,
      nios2_fpu_burst_5_upstream_readdata_from_sa => nios2_fpu_burst_5_upstream_readdata_from_sa,
      nios2_fpu_burst_5_upstream_waitrequest_from_sa => nios2_fpu_burst_5_upstream_waitrequest_from_sa,
      nios2_fpu_burst_6_upstream_readdata_from_sa => nios2_fpu_burst_6_upstream_readdata_from_sa,
      nios2_fpu_burst_6_upstream_waitrequest_from_sa => nios2_fpu_burst_6_upstream_waitrequest_from_sa,
      nios2_fpu_burst_8_upstream_readdata_from_sa => nios2_fpu_burst_8_upstream_readdata_from_sa,
      nios2_fpu_burst_8_upstream_waitrequest_from_sa => nios2_fpu_burst_8_upstream_waitrequest_from_sa,
      psw_s1_irq_from_sa => psw_s1_irq_from_sa,
      reset_n => core_clk_reset_n,
      spu_s1_irq_from_sa => spu_s1_irq_from_sa,
      systimer_s1_irq_from_sa => systimer_s1_irq_from_sa,
      sysuart_s1_irq_from_sa => sysuart_s1_irq_from_sa,
      vga_s1_irq_from_sa => vga_s1_irq_from_sa
    );


  --the_nios2_fast_fpu_instruction_master, which is an e_instance
  the_nios2_fast_fpu_instruction_master : nios2_fast_fpu_instruction_master_arbitrator
    port map(
      nios2_fast_fpu_instruction_master_address_to_slave => nios2_fast_fpu_instruction_master_address_to_slave,
      nios2_fast_fpu_instruction_master_dbs_address => nios2_fast_fpu_instruction_master_dbs_address,
      nios2_fast_fpu_instruction_master_latency_counter => nios2_fast_fpu_instruction_master_latency_counter,
      nios2_fast_fpu_instruction_master_readdata => nios2_fast_fpu_instruction_master_readdata,
      nios2_fast_fpu_instruction_master_readdatavalid => nios2_fast_fpu_instruction_master_readdatavalid,
      nios2_fast_fpu_instruction_master_waitrequest => nios2_fast_fpu_instruction_master_waitrequest,
      clk => core_clk,
      d1_nios2_fpu_burst_1_upstream_end_xfer => d1_nios2_fpu_burst_1_upstream_end_xfer,
      d1_nios2_fpu_burst_4_upstream_end_xfer => d1_nios2_fpu_burst_4_upstream_end_xfer,
      d1_nios2_fpu_burst_7_upstream_end_xfer => d1_nios2_fpu_burst_7_upstream_end_xfer,
      nios2_fast_fpu_instruction_master_address => nios2_fast_fpu_instruction_master_address,
      nios2_fast_fpu_instruction_master_burstcount => nios2_fast_fpu_instruction_master_burstcount,
      nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream => nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream,
      nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream => nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream,
      nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream => nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream,
      nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream => nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream,
      nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream => nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream,
      nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream => nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream,
      nios2_fast_fpu_instruction_master_read => nios2_fast_fpu_instruction_master_read,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register,
      nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream => nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream,
      nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream => nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream,
      nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream => nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream,
      nios2_fpu_burst_1_upstream_readdata_from_sa => nios2_fpu_burst_1_upstream_readdata_from_sa,
      nios2_fpu_burst_1_upstream_waitrequest_from_sa => nios2_fpu_burst_1_upstream_waitrequest_from_sa,
      nios2_fpu_burst_4_upstream_readdata_from_sa => nios2_fpu_burst_4_upstream_readdata_from_sa,
      nios2_fpu_burst_4_upstream_waitrequest_from_sa => nios2_fpu_burst_4_upstream_waitrequest_from_sa,
      nios2_fpu_burst_7_upstream_readdata_from_sa => nios2_fpu_burst_7_upstream_readdata_from_sa,
      nios2_fpu_burst_7_upstream_waitrequest_from_sa => nios2_fpu_burst_7_upstream_waitrequest_from_sa,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fast_fpu, which is an e_ptf_instance
  the_nios2_fast_fpu : nios2_fast_fpu
    port map(
      A_ci_multi_a => nios2_fast_fpu_custom_instruction_master_multi_a,
      A_ci_multi_b => nios2_fast_fpu_custom_instruction_master_multi_b,
      A_ci_multi_c => nios2_fast_fpu_custom_instruction_master_multi_c,
      A_ci_multi_clk_en => nios2_fast_fpu_custom_instruction_master_multi_clk_en,
      A_ci_multi_clock => nios2_fast_fpu_custom_instruction_master_multi_clk,
      A_ci_multi_dataa => nios2_fast_fpu_custom_instruction_master_multi_dataa,
      A_ci_multi_datab => nios2_fast_fpu_custom_instruction_master_multi_datab,
      A_ci_multi_estatus => nios2_fast_fpu_custom_instruction_master_multi_estatus,
      A_ci_multi_ipending => nios2_fast_fpu_custom_instruction_master_multi_ipending,
      A_ci_multi_n => nios2_fast_fpu_custom_instruction_master_multi_n,
      A_ci_multi_readra => nios2_fast_fpu_custom_instruction_master_multi_readra,
      A_ci_multi_readrb => nios2_fast_fpu_custom_instruction_master_multi_readrb,
      A_ci_multi_reset => nios2_fast_fpu_custom_instruction_master_multi_reset,
      A_ci_multi_start => nios2_fast_fpu_custom_instruction_master_multi_start,
      A_ci_multi_status => nios2_fast_fpu_custom_instruction_master_multi_status,
      A_ci_multi_writerc => nios2_fast_fpu_custom_instruction_master_multi_writerc,
      d_address => nios2_fast_fpu_data_master_address,
      d_burstcount => nios2_fast_fpu_data_master_burstcount,
      d_byteenable => nios2_fast_fpu_data_master_byteenable,
      d_read => nios2_fast_fpu_data_master_read,
      d_write => nios2_fast_fpu_data_master_write,
      d_writedata => nios2_fast_fpu_data_master_writedata,
      i_address => nios2_fast_fpu_instruction_master_address,
      i_burstcount => nios2_fast_fpu_instruction_master_burstcount,
      i_read => nios2_fast_fpu_instruction_master_read,
      jtag_debug_module_debugaccess_to_roms => nios2_fast_fpu_data_master_debugaccess,
      jtag_debug_module_readdata => nios2_fast_fpu_jtag_debug_module_readdata,
      jtag_debug_module_resetrequest => nios2_fast_fpu_jtag_debug_module_resetrequest,
      A_ci_multi_done => nios2_fast_fpu_custom_instruction_master_multi_done,
      A_ci_multi_result => nios2_fast_fpu_custom_instruction_master_multi_result,
      clk => core_clk,
      d_irq => nios2_fast_fpu_data_master_irq,
      d_readdata => nios2_fast_fpu_data_master_readdata,
      d_readdatavalid => nios2_fast_fpu_data_master_readdatavalid,
      d_waitrequest => nios2_fast_fpu_data_master_waitrequest,
      i_readdata => nios2_fast_fpu_instruction_master_readdata,
      i_readdatavalid => nios2_fast_fpu_instruction_master_readdatavalid,
      i_waitrequest => nios2_fast_fpu_instruction_master_waitrequest,
      jtag_debug_module_address => nios2_fast_fpu_jtag_debug_module_address,
      jtag_debug_module_begintransfer => nios2_fast_fpu_jtag_debug_module_begintransfer,
      jtag_debug_module_byteenable => nios2_fast_fpu_jtag_debug_module_byteenable,
      jtag_debug_module_debugaccess => nios2_fast_fpu_jtag_debug_module_debugaccess,
      jtag_debug_module_select => nios2_fast_fpu_jtag_debug_module_chipselect,
      jtag_debug_module_write => nios2_fast_fpu_jtag_debug_module_write,
      jtag_debug_module_writedata => nios2_fast_fpu_jtag_debug_module_writedata,
      reset_n => nios2_fast_fpu_custom_instruction_master_reset_n
    );


  --the_nios2_fast_fpu_fpoint_s1, which is an e_instance
  the_nios2_fast_fpu_fpoint_s1 : nios2_fast_fpu_fpoint_s1_arbitrator
    port map(
      nios2_fast_fpu_fpoint_s1_clk_en => nios2_fast_fpu_fpoint_s1_clk_en,
      nios2_fast_fpu_fpoint_s1_dataa => nios2_fast_fpu_fpoint_s1_dataa,
      nios2_fast_fpu_fpoint_s1_datab => nios2_fast_fpu_fpoint_s1_datab,
      nios2_fast_fpu_fpoint_s1_done_from_sa => nios2_fast_fpu_fpoint_s1_done_from_sa,
      nios2_fast_fpu_fpoint_s1_n => nios2_fast_fpu_fpoint_s1_n,
      nios2_fast_fpu_fpoint_s1_reset => nios2_fast_fpu_fpoint_s1_reset,
      nios2_fast_fpu_fpoint_s1_result_from_sa => nios2_fast_fpu_fpoint_s1_result_from_sa,
      nios2_fast_fpu_fpoint_s1_start => nios2_fast_fpu_fpoint_s1_start,
      clk => core_clk,
      nios2_fast_fpu_custom_instruction_master_multi_clk_en => nios2_fast_fpu_custom_instruction_master_multi_clk_en,
      nios2_fast_fpu_custom_instruction_master_multi_dataa => nios2_fast_fpu_custom_instruction_master_multi_dataa,
      nios2_fast_fpu_custom_instruction_master_multi_datab => nios2_fast_fpu_custom_instruction_master_multi_datab,
      nios2_fast_fpu_custom_instruction_master_multi_n => nios2_fast_fpu_custom_instruction_master_multi_n,
      nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_fpoint_s1 => nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_fpoint_s1,
      nios2_fast_fpu_fpoint_s1_done => nios2_fast_fpu_fpoint_s1_done,
      nios2_fast_fpu_fpoint_s1_result => nios2_fast_fpu_fpoint_s1_result,
      nios2_fast_fpu_fpoint_s1_select => nios2_fast_fpu_fpoint_s1_select,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fast_fpu_fpoint, which is an e_ptf_instance
  the_nios2_fast_fpu_fpoint : nios2_fast_fpu_fpoint
    port map(
      done => nios2_fast_fpu_fpoint_s1_done,
      result => nios2_fast_fpu_fpoint_s1_result,
      clk => core_clk,
      clk_en => nios2_fast_fpu_fpoint_s1_clk_en,
      dataa => nios2_fast_fpu_fpoint_s1_dataa,
      datab => nios2_fast_fpu_fpoint_s1_datab,
      n => nios2_fast_fpu_fpoint_s1_n,
      reset => nios2_fast_fpu_fpoint_s1_reset,
      start => nios2_fast_fpu_fpoint_s1_start
    );


  --the_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0, which is an e_instance
  the_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0 : nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_arbitrator
    port map(
      nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_clk_en => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_clk_en,
      nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_dataa => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_dataa,
      nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_datab => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_datab,
      nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done_from_sa => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done_from_sa,
      nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_n => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_n,
      nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_reset => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_reset,
      nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result_from_sa => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result_from_sa,
      nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_start => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_start,
      clk => core_clk,
      nios2_fast_fpu_custom_instruction_master_multi_clk_en => nios2_fast_fpu_custom_instruction_master_multi_clk_en,
      nios2_fast_fpu_custom_instruction_master_multi_dataa => nios2_fast_fpu_custom_instruction_master_multi_dataa,
      nios2_fast_fpu_custom_instruction_master_multi_datab => nios2_fast_fpu_custom_instruction_master_multi_datab,
      nios2_fast_fpu_custom_instruction_master_multi_n => nios2_fast_fpu_custom_instruction_master_multi_n,
      nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0 => nios2_fast_fpu_custom_instruction_master_start_nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0,
      nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done,
      nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result,
      nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_select,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fast_fpu_pixelsimd_inst, which is an e_ptf_instance
  the_nios2_fast_fpu_pixelsimd_inst : nios2_fast_fpu_pixelsimd_inst
    port map(
      done => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_done,
      result => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_result,
      clk => core_clk,
      clk_en => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_clk_en,
      dataa => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_dataa,
      datab => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_datab,
      n => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_n,
      reset => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_reset,
      start => nios2_fast_fpu_pixelsimd_inst_nios_custom_instruction_slave_0_start
    );


  --the_nios2_fpu_burst_0_upstream, which is an e_instance
  the_nios2_fpu_burst_0_upstream : nios2_fpu_burst_0_upstream_arbitrator
    port map(
      d1_nios2_fpu_burst_0_upstream_end_xfer => d1_nios2_fpu_burst_0_upstream_end_xfer,
      nios2_fpu_burst_0_upstream_address => nios2_fpu_burst_0_upstream_address,
      nios2_fpu_burst_0_upstream_burstcount => nios2_fpu_burst_0_upstream_burstcount,
      nios2_fpu_burst_0_upstream_byteaddress => nios2_fpu_burst_0_upstream_byteaddress,
      nios2_fpu_burst_0_upstream_byteenable => nios2_fpu_burst_0_upstream_byteenable,
      nios2_fpu_burst_0_upstream_debugaccess => nios2_fpu_burst_0_upstream_debugaccess,
      nios2_fpu_burst_0_upstream_read => nios2_fpu_burst_0_upstream_read,
      nios2_fpu_burst_0_upstream_readdata_from_sa => nios2_fpu_burst_0_upstream_readdata_from_sa,
      nios2_fpu_burst_0_upstream_waitrequest_from_sa => nios2_fpu_burst_0_upstream_waitrequest_from_sa,
      nios2_fpu_burst_0_upstream_write => nios2_fpu_burst_0_upstream_write,
      vga_m1_granted_nios2_fpu_burst_0_upstream => vga_m1_granted_nios2_fpu_burst_0_upstream,
      vga_m1_qualified_request_nios2_fpu_burst_0_upstream => vga_m1_qualified_request_nios2_fpu_burst_0_upstream,
      vga_m1_read_data_valid_nios2_fpu_burst_0_upstream => vga_m1_read_data_valid_nios2_fpu_burst_0_upstream,
      vga_m1_read_data_valid_nios2_fpu_burst_0_upstream_shift_register => vga_m1_read_data_valid_nios2_fpu_burst_0_upstream_shift_register,
      vga_m1_requests_nios2_fpu_burst_0_upstream => vga_m1_requests_nios2_fpu_burst_0_upstream,
      clk => core_clk,
      nios2_fpu_burst_0_upstream_readdata => nios2_fpu_burst_0_upstream_readdata,
      nios2_fpu_burst_0_upstream_readdatavalid => nios2_fpu_burst_0_upstream_readdatavalid,
      nios2_fpu_burst_0_upstream_waitrequest => nios2_fpu_burst_0_upstream_waitrequest,
      reset_n => core_clk_reset_n,
      vga_m1_address_to_slave => vga_m1_address_to_slave,
      vga_m1_burstcount => vga_m1_burstcount,
      vga_m1_dbs_address => vga_m1_dbs_address,
      vga_m1_latency_counter => vga_m1_latency_counter,
      vga_m1_read => vga_m1_read
    );


  --the_nios2_fpu_burst_0_downstream, which is an e_instance
  the_nios2_fpu_burst_0_downstream : nios2_fpu_burst_0_downstream_arbitrator
    port map(
      nios2_fpu_burst_0_downstream_address_to_slave => nios2_fpu_burst_0_downstream_address_to_slave,
      nios2_fpu_burst_0_downstream_latency_counter => nios2_fpu_burst_0_downstream_latency_counter,
      nios2_fpu_burst_0_downstream_readdata => nios2_fpu_burst_0_downstream_readdata,
      nios2_fpu_burst_0_downstream_readdatavalid => nios2_fpu_burst_0_downstream_readdatavalid,
      nios2_fpu_burst_0_downstream_reset_n => nios2_fpu_burst_0_downstream_reset_n,
      nios2_fpu_burst_0_downstream_waitrequest => nios2_fpu_burst_0_downstream_waitrequest,
      clk => core_clk,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      nios2_fpu_burst_0_downstream_address => nios2_fpu_burst_0_downstream_address,
      nios2_fpu_burst_0_downstream_burstcount => nios2_fpu_burst_0_downstream_burstcount,
      nios2_fpu_burst_0_downstream_byteenable => nios2_fpu_burst_0_downstream_byteenable,
      nios2_fpu_burst_0_downstream_granted_sdram_s1 => nios2_fpu_burst_0_downstream_granted_sdram_s1,
      nios2_fpu_burst_0_downstream_qualified_request_sdram_s1 => nios2_fpu_burst_0_downstream_qualified_request_sdram_s1,
      nios2_fpu_burst_0_downstream_read => nios2_fpu_burst_0_downstream_read,
      nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1 => nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1,
      nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1_shift_register => nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1_shift_register,
      nios2_fpu_burst_0_downstream_requests_sdram_s1 => nios2_fpu_burst_0_downstream_requests_sdram_s1,
      nios2_fpu_burst_0_downstream_write => nios2_fpu_burst_0_downstream_write,
      nios2_fpu_burst_0_downstream_writedata => nios2_fpu_burst_0_downstream_writedata,
      reset_n => core_clk_reset_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_waitrequest_from_sa => sdram_s1_waitrequest_from_sa
    );


  --the_nios2_fpu_burst_0, which is an e_ptf_instance
  the_nios2_fpu_burst_0 : nios2_fpu_burst_0
    port map(
      downstream_address => nios2_fpu_burst_0_downstream_address,
      downstream_arbitrationshare => nios2_fpu_burst_0_downstream_arbitrationshare,
      downstream_burstcount => nios2_fpu_burst_0_downstream_burstcount,
      downstream_byteenable => nios2_fpu_burst_0_downstream_byteenable,
      downstream_debugaccess => nios2_fpu_burst_0_downstream_debugaccess,
      downstream_nativeaddress => nios2_fpu_burst_0_downstream_nativeaddress,
      downstream_read => nios2_fpu_burst_0_downstream_read,
      downstream_write => nios2_fpu_burst_0_downstream_write,
      downstream_writedata => nios2_fpu_burst_0_downstream_writedata,
      upstream_readdata => nios2_fpu_burst_0_upstream_readdata,
      upstream_readdatavalid => nios2_fpu_burst_0_upstream_readdatavalid,
      upstream_waitrequest => nios2_fpu_burst_0_upstream_waitrequest,
      clk => core_clk,
      downstream_readdata => nios2_fpu_burst_0_downstream_readdata,
      downstream_readdatavalid => nios2_fpu_burst_0_downstream_readdatavalid,
      downstream_waitrequest => nios2_fpu_burst_0_downstream_waitrequest,
      reset_n => nios2_fpu_burst_0_downstream_reset_n,
      upstream_address => nios2_fpu_burst_0_upstream_byteaddress,
      upstream_burstcount => nios2_fpu_burst_0_upstream_burstcount,
      upstream_byteenable => nios2_fpu_burst_0_upstream_byteenable,
      upstream_debugaccess => nios2_fpu_burst_0_upstream_debugaccess,
      upstream_nativeaddress => nios2_fpu_burst_0_upstream_address,
      upstream_read => nios2_fpu_burst_0_upstream_read,
      upstream_write => nios2_fpu_burst_0_upstream_write,
      upstream_writedata => nios2_fpu_burst_0_upstream_writedata
    );


  --the_nios2_fpu_burst_1_upstream, which is an e_instance
  the_nios2_fpu_burst_1_upstream : nios2_fpu_burst_1_upstream_arbitrator
    port map(
      d1_nios2_fpu_burst_1_upstream_end_xfer => d1_nios2_fpu_burst_1_upstream_end_xfer,
      nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream => nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_1_upstream,
      nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream => nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_1_upstream,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register,
      nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream => nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_1_upstream,
      nios2_fpu_burst_1_upstream_address => nios2_fpu_burst_1_upstream_address,
      nios2_fpu_burst_1_upstream_byteaddress => nios2_fpu_burst_1_upstream_byteaddress,
      nios2_fpu_burst_1_upstream_byteenable => nios2_fpu_burst_1_upstream_byteenable,
      nios2_fpu_burst_1_upstream_debugaccess => nios2_fpu_burst_1_upstream_debugaccess,
      nios2_fpu_burst_1_upstream_read => nios2_fpu_burst_1_upstream_read,
      nios2_fpu_burst_1_upstream_readdata_from_sa => nios2_fpu_burst_1_upstream_readdata_from_sa,
      nios2_fpu_burst_1_upstream_waitrequest_from_sa => nios2_fpu_burst_1_upstream_waitrequest_from_sa,
      nios2_fpu_burst_1_upstream_write => nios2_fpu_burst_1_upstream_write,
      clk => core_clk,
      nios2_fast_fpu_instruction_master_address_to_slave => nios2_fast_fpu_instruction_master_address_to_slave,
      nios2_fast_fpu_instruction_master_burstcount => nios2_fast_fpu_instruction_master_burstcount,
      nios2_fast_fpu_instruction_master_dbs_address => nios2_fast_fpu_instruction_master_dbs_address,
      nios2_fast_fpu_instruction_master_latency_counter => nios2_fast_fpu_instruction_master_latency_counter,
      nios2_fast_fpu_instruction_master_read => nios2_fast_fpu_instruction_master_read,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register,
      nios2_fpu_burst_1_upstream_readdata => nios2_fpu_burst_1_upstream_readdata,
      nios2_fpu_burst_1_upstream_readdatavalid => nios2_fpu_burst_1_upstream_readdatavalid,
      nios2_fpu_burst_1_upstream_waitrequest => nios2_fpu_burst_1_upstream_waitrequest,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fpu_burst_1_downstream, which is an e_instance
  the_nios2_fpu_burst_1_downstream : nios2_fpu_burst_1_downstream_arbitrator
    port map(
      nios2_fpu_burst_1_downstream_address_to_slave => nios2_fpu_burst_1_downstream_address_to_slave,
      nios2_fpu_burst_1_downstream_latency_counter => nios2_fpu_burst_1_downstream_latency_counter,
      nios2_fpu_burst_1_downstream_readdata => nios2_fpu_burst_1_downstream_readdata,
      nios2_fpu_burst_1_downstream_readdatavalid => nios2_fpu_burst_1_downstream_readdatavalid,
      nios2_fpu_burst_1_downstream_reset_n => nios2_fpu_burst_1_downstream_reset_n,
      nios2_fpu_burst_1_downstream_waitrequest => nios2_fpu_burst_1_downstream_waitrequest,
      clk => core_clk,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      nios2_fpu_burst_1_downstream_address => nios2_fpu_burst_1_downstream_address,
      nios2_fpu_burst_1_downstream_burstcount => nios2_fpu_burst_1_downstream_burstcount,
      nios2_fpu_burst_1_downstream_byteenable => nios2_fpu_burst_1_downstream_byteenable,
      nios2_fpu_burst_1_downstream_granted_sdram_s1 => nios2_fpu_burst_1_downstream_granted_sdram_s1,
      nios2_fpu_burst_1_downstream_qualified_request_sdram_s1 => nios2_fpu_burst_1_downstream_qualified_request_sdram_s1,
      nios2_fpu_burst_1_downstream_read => nios2_fpu_burst_1_downstream_read,
      nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1 => nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1,
      nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1_shift_register => nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1_shift_register,
      nios2_fpu_burst_1_downstream_requests_sdram_s1 => nios2_fpu_burst_1_downstream_requests_sdram_s1,
      nios2_fpu_burst_1_downstream_write => nios2_fpu_burst_1_downstream_write,
      nios2_fpu_burst_1_downstream_writedata => nios2_fpu_burst_1_downstream_writedata,
      reset_n => core_clk_reset_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_waitrequest_from_sa => sdram_s1_waitrequest_from_sa
    );


  --the_nios2_fpu_burst_1, which is an e_ptf_instance
  the_nios2_fpu_burst_1 : nios2_fpu_burst_1
    port map(
      reg_downstream_address => nios2_fpu_burst_1_downstream_address,
      reg_downstream_arbitrationshare => nios2_fpu_burst_1_downstream_arbitrationshare,
      reg_downstream_burstcount => nios2_fpu_burst_1_downstream_burstcount,
      reg_downstream_byteenable => nios2_fpu_burst_1_downstream_byteenable,
      reg_downstream_debugaccess => nios2_fpu_burst_1_downstream_debugaccess,
      reg_downstream_nativeaddress => nios2_fpu_burst_1_downstream_nativeaddress,
      reg_downstream_read => nios2_fpu_burst_1_downstream_read,
      reg_downstream_write => nios2_fpu_burst_1_downstream_write,
      reg_downstream_writedata => nios2_fpu_burst_1_downstream_writedata,
      upstream_readdata => nios2_fpu_burst_1_upstream_readdata,
      upstream_readdatavalid => nios2_fpu_burst_1_upstream_readdatavalid,
      upstream_waitrequest => nios2_fpu_burst_1_upstream_waitrequest,
      clk => core_clk,
      downstream_readdata => nios2_fpu_burst_1_downstream_readdata,
      downstream_readdatavalid => nios2_fpu_burst_1_downstream_readdatavalid,
      downstream_waitrequest => nios2_fpu_burst_1_downstream_waitrequest,
      reset_n => nios2_fpu_burst_1_downstream_reset_n,
      upstream_address => nios2_fpu_burst_1_upstream_byteaddress,
      upstream_byteenable => nios2_fpu_burst_1_upstream_byteenable,
      upstream_debugaccess => nios2_fpu_burst_1_upstream_debugaccess,
      upstream_nativeaddress => nios2_fpu_burst_1_upstream_address,
      upstream_read => nios2_fpu_burst_1_upstream_read,
      upstream_write => nios2_fpu_burst_1_upstream_write,
      upstream_writedata => nios2_fpu_burst_1_upstream_writedata
    );


  --the_nios2_fpu_burst_2_upstream, which is an e_instance
  the_nios2_fpu_burst_2_upstream : nios2_fpu_burst_2_upstream_arbitrator
    port map(
      d1_nios2_fpu_burst_2_upstream_end_xfer => d1_nios2_fpu_burst_2_upstream_end_xfer,
      nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream => nios2_fast_fpu_data_master_byteenable_nios2_fpu_burst_2_upstream,
      nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream => nios2_fast_fpu_data_master_granted_nios2_fpu_burst_2_upstream,
      nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream => nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_2_upstream,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register,
      nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream => nios2_fast_fpu_data_master_requests_nios2_fpu_burst_2_upstream,
      nios2_fpu_burst_2_upstream_address => nios2_fpu_burst_2_upstream_address,
      nios2_fpu_burst_2_upstream_burstcount => nios2_fpu_burst_2_upstream_burstcount,
      nios2_fpu_burst_2_upstream_byteaddress => nios2_fpu_burst_2_upstream_byteaddress,
      nios2_fpu_burst_2_upstream_byteenable => nios2_fpu_burst_2_upstream_byteenable,
      nios2_fpu_burst_2_upstream_debugaccess => nios2_fpu_burst_2_upstream_debugaccess,
      nios2_fpu_burst_2_upstream_read => nios2_fpu_burst_2_upstream_read,
      nios2_fpu_burst_2_upstream_readdata_from_sa => nios2_fpu_burst_2_upstream_readdata_from_sa,
      nios2_fpu_burst_2_upstream_waitrequest_from_sa => nios2_fpu_burst_2_upstream_waitrequest_from_sa,
      nios2_fpu_burst_2_upstream_write => nios2_fpu_burst_2_upstream_write,
      nios2_fpu_burst_2_upstream_writedata => nios2_fpu_burst_2_upstream_writedata,
      clk => core_clk,
      nios2_fast_fpu_data_master_address_to_slave => nios2_fast_fpu_data_master_address_to_slave,
      nios2_fast_fpu_data_master_burstcount => nios2_fast_fpu_data_master_burstcount,
      nios2_fast_fpu_data_master_byteenable => nios2_fast_fpu_data_master_byteenable,
      nios2_fast_fpu_data_master_dbs_address => nios2_fast_fpu_data_master_dbs_address,
      nios2_fast_fpu_data_master_dbs_write_16 => nios2_fast_fpu_data_master_dbs_write_16,
      nios2_fast_fpu_data_master_debugaccess => nios2_fast_fpu_data_master_debugaccess,
      nios2_fast_fpu_data_master_latency_counter => nios2_fast_fpu_data_master_latency_counter,
      nios2_fast_fpu_data_master_read => nios2_fast_fpu_data_master_read,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register,
      nios2_fast_fpu_data_master_write => nios2_fast_fpu_data_master_write,
      nios2_fpu_burst_2_upstream_readdata => nios2_fpu_burst_2_upstream_readdata,
      nios2_fpu_burst_2_upstream_readdatavalid => nios2_fpu_burst_2_upstream_readdatavalid,
      nios2_fpu_burst_2_upstream_waitrequest => nios2_fpu_burst_2_upstream_waitrequest,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fpu_burst_2_downstream, which is an e_instance
  the_nios2_fpu_burst_2_downstream : nios2_fpu_burst_2_downstream_arbitrator
    port map(
      nios2_fpu_burst_2_downstream_address_to_slave => nios2_fpu_burst_2_downstream_address_to_slave,
      nios2_fpu_burst_2_downstream_latency_counter => nios2_fpu_burst_2_downstream_latency_counter,
      nios2_fpu_burst_2_downstream_readdata => nios2_fpu_burst_2_downstream_readdata,
      nios2_fpu_burst_2_downstream_readdatavalid => nios2_fpu_burst_2_downstream_readdatavalid,
      nios2_fpu_burst_2_downstream_reset_n => nios2_fpu_burst_2_downstream_reset_n,
      nios2_fpu_burst_2_downstream_waitrequest => nios2_fpu_burst_2_downstream_waitrequest,
      clk => core_clk,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      nios2_fpu_burst_2_downstream_address => nios2_fpu_burst_2_downstream_address,
      nios2_fpu_burst_2_downstream_burstcount => nios2_fpu_burst_2_downstream_burstcount,
      nios2_fpu_burst_2_downstream_byteenable => nios2_fpu_burst_2_downstream_byteenable,
      nios2_fpu_burst_2_downstream_granted_sdram_s1 => nios2_fpu_burst_2_downstream_granted_sdram_s1,
      nios2_fpu_burst_2_downstream_qualified_request_sdram_s1 => nios2_fpu_burst_2_downstream_qualified_request_sdram_s1,
      nios2_fpu_burst_2_downstream_read => nios2_fpu_burst_2_downstream_read,
      nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1 => nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1,
      nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1_shift_register => nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1_shift_register,
      nios2_fpu_burst_2_downstream_requests_sdram_s1 => nios2_fpu_burst_2_downstream_requests_sdram_s1,
      nios2_fpu_burst_2_downstream_write => nios2_fpu_burst_2_downstream_write,
      nios2_fpu_burst_2_downstream_writedata => nios2_fpu_burst_2_downstream_writedata,
      reset_n => core_clk_reset_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_waitrequest_from_sa => sdram_s1_waitrequest_from_sa
    );


  --the_nios2_fpu_burst_2, which is an e_ptf_instance
  the_nios2_fpu_burst_2 : nios2_fpu_burst_2
    port map(
      reg_downstream_address => nios2_fpu_burst_2_downstream_address,
      reg_downstream_arbitrationshare => nios2_fpu_burst_2_downstream_arbitrationshare,
      reg_downstream_burstcount => nios2_fpu_burst_2_downstream_burstcount,
      reg_downstream_byteenable => nios2_fpu_burst_2_downstream_byteenable,
      reg_downstream_debugaccess => nios2_fpu_burst_2_downstream_debugaccess,
      reg_downstream_nativeaddress => nios2_fpu_burst_2_downstream_nativeaddress,
      reg_downstream_read => nios2_fpu_burst_2_downstream_read,
      reg_downstream_write => nios2_fpu_burst_2_downstream_write,
      reg_downstream_writedata => nios2_fpu_burst_2_downstream_writedata,
      upstream_readdata => nios2_fpu_burst_2_upstream_readdata,
      upstream_readdatavalid => nios2_fpu_burst_2_upstream_readdatavalid,
      upstream_waitrequest => nios2_fpu_burst_2_upstream_waitrequest,
      clk => core_clk,
      downstream_readdata => nios2_fpu_burst_2_downstream_readdata,
      downstream_readdatavalid => nios2_fpu_burst_2_downstream_readdatavalid,
      downstream_waitrequest => nios2_fpu_burst_2_downstream_waitrequest,
      reset_n => nios2_fpu_burst_2_downstream_reset_n,
      upstream_address => nios2_fpu_burst_2_upstream_byteaddress,
      upstream_burstcount => nios2_fpu_burst_2_upstream_burstcount,
      upstream_byteenable => nios2_fpu_burst_2_upstream_byteenable,
      upstream_debugaccess => nios2_fpu_burst_2_upstream_debugaccess,
      upstream_nativeaddress => nios2_fpu_burst_2_upstream_address,
      upstream_read => nios2_fpu_burst_2_upstream_read,
      upstream_write => nios2_fpu_burst_2_upstream_write,
      upstream_writedata => nios2_fpu_burst_2_upstream_writedata
    );


  --the_nios2_fpu_burst_3_upstream, which is an e_instance
  the_nios2_fpu_burst_3_upstream : nios2_fpu_burst_3_upstream_arbitrator
    port map(
      d1_nios2_fpu_burst_3_upstream_end_xfer => d1_nios2_fpu_burst_3_upstream_end_xfer,
      nios2_fpu_burst_3_upstream_address => nios2_fpu_burst_3_upstream_address,
      nios2_fpu_burst_3_upstream_burstcount => nios2_fpu_burst_3_upstream_burstcount,
      nios2_fpu_burst_3_upstream_byteaddress => nios2_fpu_burst_3_upstream_byteaddress,
      nios2_fpu_burst_3_upstream_byteenable => nios2_fpu_burst_3_upstream_byteenable,
      nios2_fpu_burst_3_upstream_debugaccess => nios2_fpu_burst_3_upstream_debugaccess,
      nios2_fpu_burst_3_upstream_read => nios2_fpu_burst_3_upstream_read,
      nios2_fpu_burst_3_upstream_readdata_from_sa => nios2_fpu_burst_3_upstream_readdata_from_sa,
      nios2_fpu_burst_3_upstream_waitrequest_from_sa => nios2_fpu_burst_3_upstream_waitrequest_from_sa,
      nios2_fpu_burst_3_upstream_write => nios2_fpu_burst_3_upstream_write,
      spu_m1_granted_nios2_fpu_burst_3_upstream => spu_m1_granted_nios2_fpu_burst_3_upstream,
      spu_m1_qualified_request_nios2_fpu_burst_3_upstream => spu_m1_qualified_request_nios2_fpu_burst_3_upstream,
      spu_m1_read_data_valid_nios2_fpu_burst_3_upstream => spu_m1_read_data_valid_nios2_fpu_burst_3_upstream,
      spu_m1_read_data_valid_nios2_fpu_burst_3_upstream_shift_register => spu_m1_read_data_valid_nios2_fpu_burst_3_upstream_shift_register,
      spu_m1_requests_nios2_fpu_burst_3_upstream => spu_m1_requests_nios2_fpu_burst_3_upstream,
      clk => core_clk,
      nios2_fpu_burst_3_upstream_readdata => nios2_fpu_burst_3_upstream_readdata,
      nios2_fpu_burst_3_upstream_readdatavalid => nios2_fpu_burst_3_upstream_readdatavalid,
      nios2_fpu_burst_3_upstream_waitrequest => nios2_fpu_burst_3_upstream_waitrequest,
      reset_n => core_clk_reset_n,
      spu_m1_address_to_slave => spu_m1_address_to_slave,
      spu_m1_burstcount => spu_m1_burstcount,
      spu_m1_latency_counter => spu_m1_latency_counter,
      spu_m1_read => spu_m1_read
    );


  --the_nios2_fpu_burst_3_downstream, which is an e_instance
  the_nios2_fpu_burst_3_downstream : nios2_fpu_burst_3_downstream_arbitrator
    port map(
      nios2_fpu_burst_3_downstream_address_to_slave => nios2_fpu_burst_3_downstream_address_to_slave,
      nios2_fpu_burst_3_downstream_latency_counter => nios2_fpu_burst_3_downstream_latency_counter,
      nios2_fpu_burst_3_downstream_readdata => nios2_fpu_burst_3_downstream_readdata,
      nios2_fpu_burst_3_downstream_readdatavalid => nios2_fpu_burst_3_downstream_readdatavalid,
      nios2_fpu_burst_3_downstream_reset_n => nios2_fpu_burst_3_downstream_reset_n,
      nios2_fpu_burst_3_downstream_waitrequest => nios2_fpu_burst_3_downstream_waitrequest,
      clk => core_clk,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      nios2_fpu_burst_3_downstream_address => nios2_fpu_burst_3_downstream_address,
      nios2_fpu_burst_3_downstream_burstcount => nios2_fpu_burst_3_downstream_burstcount,
      nios2_fpu_burst_3_downstream_byteenable => nios2_fpu_burst_3_downstream_byteenable,
      nios2_fpu_burst_3_downstream_granted_sdram_s1 => nios2_fpu_burst_3_downstream_granted_sdram_s1,
      nios2_fpu_burst_3_downstream_qualified_request_sdram_s1 => nios2_fpu_burst_3_downstream_qualified_request_sdram_s1,
      nios2_fpu_burst_3_downstream_read => nios2_fpu_burst_3_downstream_read,
      nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1 => nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1,
      nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1_shift_register => nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1_shift_register,
      nios2_fpu_burst_3_downstream_requests_sdram_s1 => nios2_fpu_burst_3_downstream_requests_sdram_s1,
      nios2_fpu_burst_3_downstream_write => nios2_fpu_burst_3_downstream_write,
      nios2_fpu_burst_3_downstream_writedata => nios2_fpu_burst_3_downstream_writedata,
      reset_n => core_clk_reset_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_waitrequest_from_sa => sdram_s1_waitrequest_from_sa
    );


  --the_nios2_fpu_burst_3, which is an e_ptf_instance
  the_nios2_fpu_burst_3 : nios2_fpu_burst_3
    port map(
      reg_downstream_address => nios2_fpu_burst_3_downstream_address,
      reg_downstream_arbitrationshare => nios2_fpu_burst_3_downstream_arbitrationshare,
      reg_downstream_burstcount => nios2_fpu_burst_3_downstream_burstcount,
      reg_downstream_byteenable => nios2_fpu_burst_3_downstream_byteenable,
      reg_downstream_debugaccess => nios2_fpu_burst_3_downstream_debugaccess,
      reg_downstream_nativeaddress => nios2_fpu_burst_3_downstream_nativeaddress,
      reg_downstream_read => nios2_fpu_burst_3_downstream_read,
      reg_downstream_write => nios2_fpu_burst_3_downstream_write,
      reg_downstream_writedata => nios2_fpu_burst_3_downstream_writedata,
      upstream_readdata => nios2_fpu_burst_3_upstream_readdata,
      upstream_readdatavalid => nios2_fpu_burst_3_upstream_readdatavalid,
      upstream_waitrequest => nios2_fpu_burst_3_upstream_waitrequest,
      clk => core_clk,
      downstream_readdata => nios2_fpu_burst_3_downstream_readdata,
      downstream_readdatavalid => nios2_fpu_burst_3_downstream_readdatavalid,
      downstream_waitrequest => nios2_fpu_burst_3_downstream_waitrequest,
      reset_n => nios2_fpu_burst_3_downstream_reset_n,
      upstream_address => nios2_fpu_burst_3_upstream_byteaddress,
      upstream_burstcount => nios2_fpu_burst_3_upstream_burstcount,
      upstream_byteenable => nios2_fpu_burst_3_upstream_byteenable,
      upstream_debugaccess => nios2_fpu_burst_3_upstream_debugaccess,
      upstream_nativeaddress => nios2_fpu_burst_3_upstream_address,
      upstream_read => nios2_fpu_burst_3_upstream_read,
      upstream_write => nios2_fpu_burst_3_upstream_write,
      upstream_writedata => nios2_fpu_burst_3_upstream_writedata
    );


  --the_nios2_fpu_burst_4_upstream, which is an e_instance
  the_nios2_fpu_burst_4_upstream : nios2_fpu_burst_4_upstream_arbitrator
    port map(
      d1_nios2_fpu_burst_4_upstream_end_xfer => d1_nios2_fpu_burst_4_upstream_end_xfer,
      nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream => nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_4_upstream,
      nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream => nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_4_upstream,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register,
      nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream => nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_4_upstream,
      nios2_fpu_burst_4_upstream_address => nios2_fpu_burst_4_upstream_address,
      nios2_fpu_burst_4_upstream_byteaddress => nios2_fpu_burst_4_upstream_byteaddress,
      nios2_fpu_burst_4_upstream_byteenable => nios2_fpu_burst_4_upstream_byteenable,
      nios2_fpu_burst_4_upstream_debugaccess => nios2_fpu_burst_4_upstream_debugaccess,
      nios2_fpu_burst_4_upstream_read => nios2_fpu_burst_4_upstream_read,
      nios2_fpu_burst_4_upstream_readdata_from_sa => nios2_fpu_burst_4_upstream_readdata_from_sa,
      nios2_fpu_burst_4_upstream_waitrequest_from_sa => nios2_fpu_burst_4_upstream_waitrequest_from_sa,
      nios2_fpu_burst_4_upstream_write => nios2_fpu_burst_4_upstream_write,
      clk => core_clk,
      nios2_fast_fpu_instruction_master_address_to_slave => nios2_fast_fpu_instruction_master_address_to_slave,
      nios2_fast_fpu_instruction_master_burstcount => nios2_fast_fpu_instruction_master_burstcount,
      nios2_fast_fpu_instruction_master_latency_counter => nios2_fast_fpu_instruction_master_latency_counter,
      nios2_fast_fpu_instruction_master_read => nios2_fast_fpu_instruction_master_read,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register,
      nios2_fpu_burst_4_upstream_readdata => nios2_fpu_burst_4_upstream_readdata,
      nios2_fpu_burst_4_upstream_readdatavalid => nios2_fpu_burst_4_upstream_readdatavalid,
      nios2_fpu_burst_4_upstream_waitrequest => nios2_fpu_burst_4_upstream_waitrequest,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fpu_burst_4_downstream, which is an e_instance
  the_nios2_fpu_burst_4_downstream : nios2_fpu_burst_4_downstream_arbitrator
    port map(
      nios2_fpu_burst_4_downstream_address_to_slave => nios2_fpu_burst_4_downstream_address_to_slave,
      nios2_fpu_burst_4_downstream_latency_counter => nios2_fpu_burst_4_downstream_latency_counter,
      nios2_fpu_burst_4_downstream_readdata => nios2_fpu_burst_4_downstream_readdata,
      nios2_fpu_burst_4_downstream_readdatavalid => nios2_fpu_burst_4_downstream_readdatavalid,
      nios2_fpu_burst_4_downstream_reset_n => nios2_fpu_burst_4_downstream_reset_n,
      nios2_fpu_burst_4_downstream_waitrequest => nios2_fpu_burst_4_downstream_waitrequest,
      clk => core_clk,
      d1_nios2_fast_fpu_jtag_debug_module_end_xfer => d1_nios2_fast_fpu_jtag_debug_module_end_xfer,
      nios2_fast_fpu_jtag_debug_module_readdata_from_sa => nios2_fast_fpu_jtag_debug_module_readdata_from_sa,
      nios2_fpu_burst_4_downstream_address => nios2_fpu_burst_4_downstream_address,
      nios2_fpu_burst_4_downstream_burstcount => nios2_fpu_burst_4_downstream_burstcount,
      nios2_fpu_burst_4_downstream_byteenable => nios2_fpu_burst_4_downstream_byteenable,
      nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_4_downstream_granted_nios2_fast_fpu_jtag_debug_module,
      nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_4_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module,
      nios2_fpu_burst_4_downstream_read => nios2_fpu_burst_4_downstream_read,
      nios2_fpu_burst_4_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_4_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module,
      nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_4_downstream_requests_nios2_fast_fpu_jtag_debug_module,
      nios2_fpu_burst_4_downstream_write => nios2_fpu_burst_4_downstream_write,
      nios2_fpu_burst_4_downstream_writedata => nios2_fpu_burst_4_downstream_writedata,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fpu_burst_4, which is an e_ptf_instance
  the_nios2_fpu_burst_4 : nios2_fpu_burst_4
    port map(
      reg_downstream_address => nios2_fpu_burst_4_downstream_address,
      reg_downstream_arbitrationshare => nios2_fpu_burst_4_downstream_arbitrationshare,
      reg_downstream_burstcount => nios2_fpu_burst_4_downstream_burstcount,
      reg_downstream_byteenable => nios2_fpu_burst_4_downstream_byteenable,
      reg_downstream_debugaccess => nios2_fpu_burst_4_downstream_debugaccess,
      reg_downstream_nativeaddress => nios2_fpu_burst_4_downstream_nativeaddress,
      reg_downstream_read => nios2_fpu_burst_4_downstream_read,
      reg_downstream_write => nios2_fpu_burst_4_downstream_write,
      reg_downstream_writedata => nios2_fpu_burst_4_downstream_writedata,
      upstream_readdata => nios2_fpu_burst_4_upstream_readdata,
      upstream_readdatavalid => nios2_fpu_burst_4_upstream_readdatavalid,
      upstream_waitrequest => nios2_fpu_burst_4_upstream_waitrequest,
      clk => core_clk,
      downstream_readdata => nios2_fpu_burst_4_downstream_readdata,
      downstream_readdatavalid => nios2_fpu_burst_4_downstream_readdatavalid,
      downstream_waitrequest => nios2_fpu_burst_4_downstream_waitrequest,
      reset_n => nios2_fpu_burst_4_downstream_reset_n,
      upstream_address => nios2_fpu_burst_4_upstream_byteaddress,
      upstream_byteenable => nios2_fpu_burst_4_upstream_byteenable,
      upstream_debugaccess => nios2_fpu_burst_4_upstream_debugaccess,
      upstream_nativeaddress => nios2_fpu_burst_4_upstream_address,
      upstream_read => nios2_fpu_burst_4_upstream_read,
      upstream_write => nios2_fpu_burst_4_upstream_write,
      upstream_writedata => nios2_fpu_burst_4_upstream_writedata
    );


  --the_nios2_fpu_burst_5_upstream, which is an e_instance
  the_nios2_fpu_burst_5_upstream : nios2_fpu_burst_5_upstream_arbitrator
    port map(
      d1_nios2_fpu_burst_5_upstream_end_xfer => d1_nios2_fpu_burst_5_upstream_end_xfer,
      nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream => nios2_fast_fpu_data_master_granted_nios2_fpu_burst_5_upstream,
      nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream => nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_5_upstream,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register,
      nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream => nios2_fast_fpu_data_master_requests_nios2_fpu_burst_5_upstream,
      nios2_fpu_burst_5_upstream_address => nios2_fpu_burst_5_upstream_address,
      nios2_fpu_burst_5_upstream_burstcount => nios2_fpu_burst_5_upstream_burstcount,
      nios2_fpu_burst_5_upstream_byteaddress => nios2_fpu_burst_5_upstream_byteaddress,
      nios2_fpu_burst_5_upstream_byteenable => nios2_fpu_burst_5_upstream_byteenable,
      nios2_fpu_burst_5_upstream_debugaccess => nios2_fpu_burst_5_upstream_debugaccess,
      nios2_fpu_burst_5_upstream_read => nios2_fpu_burst_5_upstream_read,
      nios2_fpu_burst_5_upstream_readdata_from_sa => nios2_fpu_burst_5_upstream_readdata_from_sa,
      nios2_fpu_burst_5_upstream_waitrequest_from_sa => nios2_fpu_burst_5_upstream_waitrequest_from_sa,
      nios2_fpu_burst_5_upstream_write => nios2_fpu_burst_5_upstream_write,
      nios2_fpu_burst_5_upstream_writedata => nios2_fpu_burst_5_upstream_writedata,
      clk => core_clk,
      nios2_fast_fpu_data_master_address_to_slave => nios2_fast_fpu_data_master_address_to_slave,
      nios2_fast_fpu_data_master_burstcount => nios2_fast_fpu_data_master_burstcount,
      nios2_fast_fpu_data_master_byteenable => nios2_fast_fpu_data_master_byteenable,
      nios2_fast_fpu_data_master_debugaccess => nios2_fast_fpu_data_master_debugaccess,
      nios2_fast_fpu_data_master_latency_counter => nios2_fast_fpu_data_master_latency_counter,
      nios2_fast_fpu_data_master_read => nios2_fast_fpu_data_master_read,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register,
      nios2_fast_fpu_data_master_write => nios2_fast_fpu_data_master_write,
      nios2_fast_fpu_data_master_writedata => nios2_fast_fpu_data_master_writedata,
      nios2_fpu_burst_5_upstream_readdata => nios2_fpu_burst_5_upstream_readdata,
      nios2_fpu_burst_5_upstream_readdatavalid => nios2_fpu_burst_5_upstream_readdatavalid,
      nios2_fpu_burst_5_upstream_waitrequest => nios2_fpu_burst_5_upstream_waitrequest,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fpu_burst_5_downstream, which is an e_instance
  the_nios2_fpu_burst_5_downstream : nios2_fpu_burst_5_downstream_arbitrator
    port map(
      nios2_fpu_burst_5_downstream_address_to_slave => nios2_fpu_burst_5_downstream_address_to_slave,
      nios2_fpu_burst_5_downstream_latency_counter => nios2_fpu_burst_5_downstream_latency_counter,
      nios2_fpu_burst_5_downstream_readdata => nios2_fpu_burst_5_downstream_readdata,
      nios2_fpu_burst_5_downstream_readdatavalid => nios2_fpu_burst_5_downstream_readdatavalid,
      nios2_fpu_burst_5_downstream_reset_n => nios2_fpu_burst_5_downstream_reset_n,
      nios2_fpu_burst_5_downstream_waitrequest => nios2_fpu_burst_5_downstream_waitrequest,
      clk => core_clk,
      d1_nios2_fast_fpu_jtag_debug_module_end_xfer => d1_nios2_fast_fpu_jtag_debug_module_end_xfer,
      nios2_fast_fpu_jtag_debug_module_readdata_from_sa => nios2_fast_fpu_jtag_debug_module_readdata_from_sa,
      nios2_fpu_burst_5_downstream_address => nios2_fpu_burst_5_downstream_address,
      nios2_fpu_burst_5_downstream_burstcount => nios2_fpu_burst_5_downstream_burstcount,
      nios2_fpu_burst_5_downstream_byteenable => nios2_fpu_burst_5_downstream_byteenable,
      nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_5_downstream_granted_nios2_fast_fpu_jtag_debug_module,
      nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_5_downstream_qualified_request_nios2_fast_fpu_jtag_debug_module,
      nios2_fpu_burst_5_downstream_read => nios2_fpu_burst_5_downstream_read,
      nios2_fpu_burst_5_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_5_downstream_read_data_valid_nios2_fast_fpu_jtag_debug_module,
      nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module => nios2_fpu_burst_5_downstream_requests_nios2_fast_fpu_jtag_debug_module,
      nios2_fpu_burst_5_downstream_write => nios2_fpu_burst_5_downstream_write,
      nios2_fpu_burst_5_downstream_writedata => nios2_fpu_burst_5_downstream_writedata,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fpu_burst_5, which is an e_ptf_instance
  the_nios2_fpu_burst_5 : nios2_fpu_burst_5
    port map(
      reg_downstream_address => nios2_fpu_burst_5_downstream_address,
      reg_downstream_arbitrationshare => nios2_fpu_burst_5_downstream_arbitrationshare,
      reg_downstream_burstcount => nios2_fpu_burst_5_downstream_burstcount,
      reg_downstream_byteenable => nios2_fpu_burst_5_downstream_byteenable,
      reg_downstream_debugaccess => nios2_fpu_burst_5_downstream_debugaccess,
      reg_downstream_nativeaddress => nios2_fpu_burst_5_downstream_nativeaddress,
      reg_downstream_read => nios2_fpu_burst_5_downstream_read,
      reg_downstream_write => nios2_fpu_burst_5_downstream_write,
      reg_downstream_writedata => nios2_fpu_burst_5_downstream_writedata,
      upstream_readdata => nios2_fpu_burst_5_upstream_readdata,
      upstream_readdatavalid => nios2_fpu_burst_5_upstream_readdatavalid,
      upstream_waitrequest => nios2_fpu_burst_5_upstream_waitrequest,
      clk => core_clk,
      downstream_readdata => nios2_fpu_burst_5_downstream_readdata,
      downstream_readdatavalid => nios2_fpu_burst_5_downstream_readdatavalid,
      downstream_waitrequest => nios2_fpu_burst_5_downstream_waitrequest,
      reset_n => nios2_fpu_burst_5_downstream_reset_n,
      upstream_address => nios2_fpu_burst_5_upstream_byteaddress,
      upstream_burstcount => nios2_fpu_burst_5_upstream_burstcount,
      upstream_byteenable => nios2_fpu_burst_5_upstream_byteenable,
      upstream_debugaccess => nios2_fpu_burst_5_upstream_debugaccess,
      upstream_nativeaddress => nios2_fpu_burst_5_upstream_address,
      upstream_read => nios2_fpu_burst_5_upstream_read,
      upstream_write => nios2_fpu_burst_5_upstream_write,
      upstream_writedata => nios2_fpu_burst_5_upstream_writedata
    );


  --the_nios2_fpu_burst_6_upstream, which is an e_instance
  the_nios2_fpu_burst_6_upstream : nios2_fpu_burst_6_upstream_arbitrator
    port map(
      d1_nios2_fpu_burst_6_upstream_end_xfer => d1_nios2_fpu_burst_6_upstream_end_xfer,
      nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream => nios2_fast_fpu_data_master_granted_nios2_fpu_burst_6_upstream,
      nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream => nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_6_upstream,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register,
      nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream => nios2_fast_fpu_data_master_requests_nios2_fpu_burst_6_upstream,
      nios2_fpu_burst_6_upstream_address => nios2_fpu_burst_6_upstream_address,
      nios2_fpu_burst_6_upstream_burstcount => nios2_fpu_burst_6_upstream_burstcount,
      nios2_fpu_burst_6_upstream_byteaddress => nios2_fpu_burst_6_upstream_byteaddress,
      nios2_fpu_burst_6_upstream_byteenable => nios2_fpu_burst_6_upstream_byteenable,
      nios2_fpu_burst_6_upstream_debugaccess => nios2_fpu_burst_6_upstream_debugaccess,
      nios2_fpu_burst_6_upstream_read => nios2_fpu_burst_6_upstream_read,
      nios2_fpu_burst_6_upstream_readdata_from_sa => nios2_fpu_burst_6_upstream_readdata_from_sa,
      nios2_fpu_burst_6_upstream_waitrequest_from_sa => nios2_fpu_burst_6_upstream_waitrequest_from_sa,
      nios2_fpu_burst_6_upstream_write => nios2_fpu_burst_6_upstream_write,
      nios2_fpu_burst_6_upstream_writedata => nios2_fpu_burst_6_upstream_writedata,
      clk => core_clk,
      nios2_fast_fpu_data_master_address_to_slave => nios2_fast_fpu_data_master_address_to_slave,
      nios2_fast_fpu_data_master_burstcount => nios2_fast_fpu_data_master_burstcount,
      nios2_fast_fpu_data_master_byteenable => nios2_fast_fpu_data_master_byteenable,
      nios2_fast_fpu_data_master_debugaccess => nios2_fast_fpu_data_master_debugaccess,
      nios2_fast_fpu_data_master_latency_counter => nios2_fast_fpu_data_master_latency_counter,
      nios2_fast_fpu_data_master_read => nios2_fast_fpu_data_master_read,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register,
      nios2_fast_fpu_data_master_write => nios2_fast_fpu_data_master_write,
      nios2_fast_fpu_data_master_writedata => nios2_fast_fpu_data_master_writedata,
      nios2_fpu_burst_6_upstream_readdata => nios2_fpu_burst_6_upstream_readdata,
      nios2_fpu_burst_6_upstream_readdatavalid => nios2_fpu_burst_6_upstream_readdatavalid,
      nios2_fpu_burst_6_upstream_waitrequest => nios2_fpu_burst_6_upstream_waitrequest,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fpu_burst_6_downstream, which is an e_instance
  the_nios2_fpu_burst_6_downstream : nios2_fpu_burst_6_downstream_arbitrator
    port map(
      nios2_fpu_burst_6_downstream_address_to_slave => nios2_fpu_burst_6_downstream_address_to_slave,
      nios2_fpu_burst_6_downstream_latency_counter => nios2_fpu_burst_6_downstream_latency_counter,
      nios2_fpu_burst_6_downstream_readdata => nios2_fpu_burst_6_downstream_readdata,
      nios2_fpu_burst_6_downstream_readdatavalid => nios2_fpu_burst_6_downstream_readdatavalid,
      nios2_fpu_burst_6_downstream_reset_n => nios2_fpu_burst_6_downstream_reset_n,
      nios2_fpu_burst_6_downstream_waitrequest => nios2_fpu_burst_6_downstream_waitrequest,
      clk => core_clk,
      d1_ipl_memory_s1_end_xfer => d1_ipl_memory_s1_end_xfer,
      ipl_memory_s1_readdata_from_sa => ipl_memory_s1_readdata_from_sa,
      nios2_fpu_burst_6_downstream_address => nios2_fpu_burst_6_downstream_address,
      nios2_fpu_burst_6_downstream_burstcount => nios2_fpu_burst_6_downstream_burstcount,
      nios2_fpu_burst_6_downstream_byteenable => nios2_fpu_burst_6_downstream_byteenable,
      nios2_fpu_burst_6_downstream_granted_ipl_memory_s1 => nios2_fpu_burst_6_downstream_granted_ipl_memory_s1,
      nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1 => nios2_fpu_burst_6_downstream_qualified_request_ipl_memory_s1,
      nios2_fpu_burst_6_downstream_read => nios2_fpu_burst_6_downstream_read,
      nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1 => nios2_fpu_burst_6_downstream_read_data_valid_ipl_memory_s1,
      nios2_fpu_burst_6_downstream_requests_ipl_memory_s1 => nios2_fpu_burst_6_downstream_requests_ipl_memory_s1,
      nios2_fpu_burst_6_downstream_write => nios2_fpu_burst_6_downstream_write,
      nios2_fpu_burst_6_downstream_writedata => nios2_fpu_burst_6_downstream_writedata,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fpu_burst_6, which is an e_ptf_instance
  the_nios2_fpu_burst_6 : nios2_fpu_burst_6
    port map(
      reg_downstream_address => nios2_fpu_burst_6_downstream_address,
      reg_downstream_arbitrationshare => nios2_fpu_burst_6_downstream_arbitrationshare,
      reg_downstream_burstcount => nios2_fpu_burst_6_downstream_burstcount,
      reg_downstream_byteenable => nios2_fpu_burst_6_downstream_byteenable,
      reg_downstream_debugaccess => nios2_fpu_burst_6_downstream_debugaccess,
      reg_downstream_nativeaddress => nios2_fpu_burst_6_downstream_nativeaddress,
      reg_downstream_read => nios2_fpu_burst_6_downstream_read,
      reg_downstream_write => nios2_fpu_burst_6_downstream_write,
      reg_downstream_writedata => nios2_fpu_burst_6_downstream_writedata,
      upstream_readdata => nios2_fpu_burst_6_upstream_readdata,
      upstream_readdatavalid => nios2_fpu_burst_6_upstream_readdatavalid,
      upstream_waitrequest => nios2_fpu_burst_6_upstream_waitrequest,
      clk => core_clk,
      downstream_readdata => nios2_fpu_burst_6_downstream_readdata,
      downstream_readdatavalid => nios2_fpu_burst_6_downstream_readdatavalid,
      downstream_waitrequest => nios2_fpu_burst_6_downstream_waitrequest,
      reset_n => nios2_fpu_burst_6_downstream_reset_n,
      upstream_address => nios2_fpu_burst_6_upstream_byteaddress,
      upstream_burstcount => nios2_fpu_burst_6_upstream_burstcount,
      upstream_byteenable => nios2_fpu_burst_6_upstream_byteenable,
      upstream_debugaccess => nios2_fpu_burst_6_upstream_debugaccess,
      upstream_nativeaddress => nios2_fpu_burst_6_upstream_address,
      upstream_read => nios2_fpu_burst_6_upstream_read,
      upstream_write => nios2_fpu_burst_6_upstream_write,
      upstream_writedata => nios2_fpu_burst_6_upstream_writedata
    );


  --the_nios2_fpu_burst_7_upstream, which is an e_instance
  the_nios2_fpu_burst_7_upstream : nios2_fpu_burst_7_upstream_arbitrator
    port map(
      d1_nios2_fpu_burst_7_upstream_end_xfer => d1_nios2_fpu_burst_7_upstream_end_xfer,
      nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream => nios2_fast_fpu_instruction_master_granted_nios2_fpu_burst_7_upstream,
      nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream => nios2_fast_fpu_instruction_master_qualified_request_nios2_fpu_burst_7_upstream,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_7_upstream_shift_register,
      nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream => nios2_fast_fpu_instruction_master_requests_nios2_fpu_burst_7_upstream,
      nios2_fpu_burst_7_upstream_address => nios2_fpu_burst_7_upstream_address,
      nios2_fpu_burst_7_upstream_byteaddress => nios2_fpu_burst_7_upstream_byteaddress,
      nios2_fpu_burst_7_upstream_byteenable => nios2_fpu_burst_7_upstream_byteenable,
      nios2_fpu_burst_7_upstream_debugaccess => nios2_fpu_burst_7_upstream_debugaccess,
      nios2_fpu_burst_7_upstream_read => nios2_fpu_burst_7_upstream_read,
      nios2_fpu_burst_7_upstream_readdata_from_sa => nios2_fpu_burst_7_upstream_readdata_from_sa,
      nios2_fpu_burst_7_upstream_waitrequest_from_sa => nios2_fpu_burst_7_upstream_waitrequest_from_sa,
      nios2_fpu_burst_7_upstream_write => nios2_fpu_burst_7_upstream_write,
      clk => core_clk,
      nios2_fast_fpu_instruction_master_address_to_slave => nios2_fast_fpu_instruction_master_address_to_slave,
      nios2_fast_fpu_instruction_master_burstcount => nios2_fast_fpu_instruction_master_burstcount,
      nios2_fast_fpu_instruction_master_latency_counter => nios2_fast_fpu_instruction_master_latency_counter,
      nios2_fast_fpu_instruction_master_read => nios2_fast_fpu_instruction_master_read,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_1_upstream_shift_register,
      nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register => nios2_fast_fpu_instruction_master_read_data_valid_nios2_fpu_burst_4_upstream_shift_register,
      nios2_fpu_burst_7_upstream_readdata => nios2_fpu_burst_7_upstream_readdata,
      nios2_fpu_burst_7_upstream_readdatavalid => nios2_fpu_burst_7_upstream_readdatavalid,
      nios2_fpu_burst_7_upstream_waitrequest => nios2_fpu_burst_7_upstream_waitrequest,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fpu_burst_7_downstream, which is an e_instance
  the_nios2_fpu_burst_7_downstream : nios2_fpu_burst_7_downstream_arbitrator
    port map(
      nios2_fpu_burst_7_downstream_address_to_slave => nios2_fpu_burst_7_downstream_address_to_slave,
      nios2_fpu_burst_7_downstream_latency_counter => nios2_fpu_burst_7_downstream_latency_counter,
      nios2_fpu_burst_7_downstream_readdata => nios2_fpu_burst_7_downstream_readdata,
      nios2_fpu_burst_7_downstream_readdatavalid => nios2_fpu_burst_7_downstream_readdatavalid,
      nios2_fpu_burst_7_downstream_reset_n => nios2_fpu_burst_7_downstream_reset_n,
      nios2_fpu_burst_7_downstream_waitrequest => nios2_fpu_burst_7_downstream_waitrequest,
      clk => core_clk,
      d1_ipl_memory_s1_end_xfer => d1_ipl_memory_s1_end_xfer,
      ipl_memory_s1_readdata_from_sa => ipl_memory_s1_readdata_from_sa,
      nios2_fpu_burst_7_downstream_address => nios2_fpu_burst_7_downstream_address,
      nios2_fpu_burst_7_downstream_burstcount => nios2_fpu_burst_7_downstream_burstcount,
      nios2_fpu_burst_7_downstream_byteenable => nios2_fpu_burst_7_downstream_byteenable,
      nios2_fpu_burst_7_downstream_granted_ipl_memory_s1 => nios2_fpu_burst_7_downstream_granted_ipl_memory_s1,
      nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1 => nios2_fpu_burst_7_downstream_qualified_request_ipl_memory_s1,
      nios2_fpu_burst_7_downstream_read => nios2_fpu_burst_7_downstream_read,
      nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1 => nios2_fpu_burst_7_downstream_read_data_valid_ipl_memory_s1,
      nios2_fpu_burst_7_downstream_requests_ipl_memory_s1 => nios2_fpu_burst_7_downstream_requests_ipl_memory_s1,
      nios2_fpu_burst_7_downstream_write => nios2_fpu_burst_7_downstream_write,
      nios2_fpu_burst_7_downstream_writedata => nios2_fpu_burst_7_downstream_writedata,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fpu_burst_7, which is an e_ptf_instance
  the_nios2_fpu_burst_7 : nios2_fpu_burst_7
    port map(
      reg_downstream_address => nios2_fpu_burst_7_downstream_address,
      reg_downstream_arbitrationshare => nios2_fpu_burst_7_downstream_arbitrationshare,
      reg_downstream_burstcount => nios2_fpu_burst_7_downstream_burstcount,
      reg_downstream_byteenable => nios2_fpu_burst_7_downstream_byteenable,
      reg_downstream_debugaccess => nios2_fpu_burst_7_downstream_debugaccess,
      reg_downstream_nativeaddress => nios2_fpu_burst_7_downstream_nativeaddress,
      reg_downstream_read => nios2_fpu_burst_7_downstream_read,
      reg_downstream_write => nios2_fpu_burst_7_downstream_write,
      reg_downstream_writedata => nios2_fpu_burst_7_downstream_writedata,
      upstream_readdata => nios2_fpu_burst_7_upstream_readdata,
      upstream_readdatavalid => nios2_fpu_burst_7_upstream_readdatavalid,
      upstream_waitrequest => nios2_fpu_burst_7_upstream_waitrequest,
      clk => core_clk,
      downstream_readdata => nios2_fpu_burst_7_downstream_readdata,
      downstream_readdatavalid => nios2_fpu_burst_7_downstream_readdatavalid,
      downstream_waitrequest => nios2_fpu_burst_7_downstream_waitrequest,
      reset_n => nios2_fpu_burst_7_downstream_reset_n,
      upstream_address => nios2_fpu_burst_7_upstream_byteaddress,
      upstream_byteenable => nios2_fpu_burst_7_upstream_byteenable,
      upstream_debugaccess => nios2_fpu_burst_7_upstream_debugaccess,
      upstream_nativeaddress => nios2_fpu_burst_7_upstream_address,
      upstream_read => nios2_fpu_burst_7_upstream_read,
      upstream_write => nios2_fpu_burst_7_upstream_write,
      upstream_writedata => nios2_fpu_burst_7_upstream_writedata
    );


  --the_nios2_fpu_burst_8_upstream, which is an e_instance
  the_nios2_fpu_burst_8_upstream : nios2_fpu_burst_8_upstream_arbitrator
    port map(
      d1_nios2_fpu_burst_8_upstream_end_xfer => d1_nios2_fpu_burst_8_upstream_end_xfer,
      nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream => nios2_fast_fpu_data_master_granted_nios2_fpu_burst_8_upstream,
      nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream => nios2_fast_fpu_data_master_qualified_request_nios2_fpu_burst_8_upstream,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_8_upstream_shift_register,
      nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream => nios2_fast_fpu_data_master_requests_nios2_fpu_burst_8_upstream,
      nios2_fpu_burst_8_upstream_address => nios2_fpu_burst_8_upstream_address,
      nios2_fpu_burst_8_upstream_burstcount => nios2_fpu_burst_8_upstream_burstcount,
      nios2_fpu_burst_8_upstream_byteaddress => nios2_fpu_burst_8_upstream_byteaddress,
      nios2_fpu_burst_8_upstream_byteenable => nios2_fpu_burst_8_upstream_byteenable,
      nios2_fpu_burst_8_upstream_debugaccess => nios2_fpu_burst_8_upstream_debugaccess,
      nios2_fpu_burst_8_upstream_read => nios2_fpu_burst_8_upstream_read,
      nios2_fpu_burst_8_upstream_readdata_from_sa => nios2_fpu_burst_8_upstream_readdata_from_sa,
      nios2_fpu_burst_8_upstream_waitrequest_from_sa => nios2_fpu_burst_8_upstream_waitrequest_from_sa,
      nios2_fpu_burst_8_upstream_write => nios2_fpu_burst_8_upstream_write,
      nios2_fpu_burst_8_upstream_writedata => nios2_fpu_burst_8_upstream_writedata,
      clk => core_clk,
      nios2_fast_fpu_data_master_address_to_slave => nios2_fast_fpu_data_master_address_to_slave,
      nios2_fast_fpu_data_master_burstcount => nios2_fast_fpu_data_master_burstcount,
      nios2_fast_fpu_data_master_byteenable => nios2_fast_fpu_data_master_byteenable,
      nios2_fast_fpu_data_master_debugaccess => nios2_fast_fpu_data_master_debugaccess,
      nios2_fast_fpu_data_master_latency_counter => nios2_fast_fpu_data_master_latency_counter,
      nios2_fast_fpu_data_master_read => nios2_fast_fpu_data_master_read,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_2_upstream_shift_register,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_5_upstream_shift_register,
      nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register => nios2_fast_fpu_data_master_read_data_valid_nios2_fpu_burst_6_upstream_shift_register,
      nios2_fast_fpu_data_master_write => nios2_fast_fpu_data_master_write,
      nios2_fast_fpu_data_master_writedata => nios2_fast_fpu_data_master_writedata,
      nios2_fpu_burst_8_upstream_readdata => nios2_fpu_burst_8_upstream_readdata,
      nios2_fpu_burst_8_upstream_readdatavalid => nios2_fpu_burst_8_upstream_readdatavalid,
      nios2_fpu_burst_8_upstream_waitrequest => nios2_fpu_burst_8_upstream_waitrequest,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fpu_burst_8_downstream, which is an e_instance
  the_nios2_fpu_burst_8_downstream : nios2_fpu_burst_8_downstream_arbitrator
    port map(
      nios2_fpu_burst_8_downstream_address_to_slave => nios2_fpu_burst_8_downstream_address_to_slave,
      nios2_fpu_burst_8_downstream_latency_counter => nios2_fpu_burst_8_downstream_latency_counter,
      nios2_fpu_burst_8_downstream_readdata => nios2_fpu_burst_8_downstream_readdata,
      nios2_fpu_burst_8_downstream_readdatavalid => nios2_fpu_burst_8_downstream_readdatavalid,
      nios2_fpu_burst_8_downstream_reset_n => nios2_fpu_burst_8_downstream_reset_n,
      nios2_fpu_burst_8_downstream_waitrequest => nios2_fpu_burst_8_downstream_waitrequest,
      clk => core_clk,
      d1_nios2_fpu_clock_0_in_end_xfer => d1_nios2_fpu_clock_0_in_end_xfer,
      nios2_fpu_burst_8_downstream_address => nios2_fpu_burst_8_downstream_address,
      nios2_fpu_burst_8_downstream_burstcount => nios2_fpu_burst_8_downstream_burstcount,
      nios2_fpu_burst_8_downstream_byteenable => nios2_fpu_burst_8_downstream_byteenable,
      nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in => nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in,
      nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in => nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in,
      nios2_fpu_burst_8_downstream_read => nios2_fpu_burst_8_downstream_read,
      nios2_fpu_burst_8_downstream_read_data_valid_nios2_fpu_clock_0_in => nios2_fpu_burst_8_downstream_read_data_valid_nios2_fpu_clock_0_in,
      nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in => nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in,
      nios2_fpu_burst_8_downstream_write => nios2_fpu_burst_8_downstream_write,
      nios2_fpu_burst_8_downstream_writedata => nios2_fpu_burst_8_downstream_writedata,
      nios2_fpu_clock_0_in_readdata_from_sa => nios2_fpu_clock_0_in_readdata_from_sa,
      nios2_fpu_clock_0_in_waitrequest_from_sa => nios2_fpu_clock_0_in_waitrequest_from_sa,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fpu_burst_8, which is an e_ptf_instance
  the_nios2_fpu_burst_8 : nios2_fpu_burst_8
    port map(
      reg_downstream_address => nios2_fpu_burst_8_downstream_address,
      reg_downstream_arbitrationshare => nios2_fpu_burst_8_downstream_arbitrationshare,
      reg_downstream_burstcount => nios2_fpu_burst_8_downstream_burstcount,
      reg_downstream_byteenable => nios2_fpu_burst_8_downstream_byteenable,
      reg_downstream_debugaccess => nios2_fpu_burst_8_downstream_debugaccess,
      reg_downstream_nativeaddress => nios2_fpu_burst_8_downstream_nativeaddress,
      reg_downstream_read => nios2_fpu_burst_8_downstream_read,
      reg_downstream_write => nios2_fpu_burst_8_downstream_write,
      reg_downstream_writedata => nios2_fpu_burst_8_downstream_writedata,
      upstream_readdata => nios2_fpu_burst_8_upstream_readdata,
      upstream_readdatavalid => nios2_fpu_burst_8_upstream_readdatavalid,
      upstream_waitrequest => nios2_fpu_burst_8_upstream_waitrequest,
      clk => core_clk,
      downstream_readdata => nios2_fpu_burst_8_downstream_readdata,
      downstream_readdatavalid => nios2_fpu_burst_8_downstream_readdatavalid,
      downstream_waitrequest => nios2_fpu_burst_8_downstream_waitrequest,
      reset_n => nios2_fpu_burst_8_downstream_reset_n,
      upstream_address => nios2_fpu_burst_8_upstream_byteaddress,
      upstream_burstcount => nios2_fpu_burst_8_upstream_burstcount,
      upstream_byteenable => nios2_fpu_burst_8_upstream_byteenable,
      upstream_debugaccess => nios2_fpu_burst_8_upstream_debugaccess,
      upstream_nativeaddress => nios2_fpu_burst_8_upstream_address,
      upstream_read => nios2_fpu_burst_8_upstream_read,
      upstream_write => nios2_fpu_burst_8_upstream_write,
      upstream_writedata => nios2_fpu_burst_8_upstream_writedata
    );


  --the_nios2_fpu_clock_0_in, which is an e_instance
  the_nios2_fpu_clock_0_in : nios2_fpu_clock_0_in_arbitrator
    port map(
      d1_nios2_fpu_clock_0_in_end_xfer => d1_nios2_fpu_clock_0_in_end_xfer,
      nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in => nios2_fpu_burst_8_downstream_granted_nios2_fpu_clock_0_in,
      nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in => nios2_fpu_burst_8_downstream_qualified_request_nios2_fpu_clock_0_in,
      nios2_fpu_burst_8_downstream_read_data_valid_nios2_fpu_clock_0_in => nios2_fpu_burst_8_downstream_read_data_valid_nios2_fpu_clock_0_in,
      nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in => nios2_fpu_burst_8_downstream_requests_nios2_fpu_clock_0_in,
      nios2_fpu_clock_0_in_address => nios2_fpu_clock_0_in_address,
      nios2_fpu_clock_0_in_byteenable => nios2_fpu_clock_0_in_byteenable,
      nios2_fpu_clock_0_in_endofpacket_from_sa => nios2_fpu_clock_0_in_endofpacket_from_sa,
      nios2_fpu_clock_0_in_nativeaddress => nios2_fpu_clock_0_in_nativeaddress,
      nios2_fpu_clock_0_in_read => nios2_fpu_clock_0_in_read,
      nios2_fpu_clock_0_in_readdata_from_sa => nios2_fpu_clock_0_in_readdata_from_sa,
      nios2_fpu_clock_0_in_reset_n => nios2_fpu_clock_0_in_reset_n,
      nios2_fpu_clock_0_in_waitrequest_from_sa => nios2_fpu_clock_0_in_waitrequest_from_sa,
      nios2_fpu_clock_0_in_write => nios2_fpu_clock_0_in_write,
      nios2_fpu_clock_0_in_writedata => nios2_fpu_clock_0_in_writedata,
      clk => core_clk,
      nios2_fpu_burst_8_downstream_address_to_slave => nios2_fpu_burst_8_downstream_address_to_slave,
      nios2_fpu_burst_8_downstream_arbitrationshare => nios2_fpu_burst_8_downstream_arbitrationshare,
      nios2_fpu_burst_8_downstream_burstcount => nios2_fpu_burst_8_downstream_burstcount,
      nios2_fpu_burst_8_downstream_byteenable => nios2_fpu_burst_8_downstream_byteenable,
      nios2_fpu_burst_8_downstream_latency_counter => nios2_fpu_burst_8_downstream_latency_counter,
      nios2_fpu_burst_8_downstream_nativeaddress => nios2_fpu_burst_8_downstream_nativeaddress,
      nios2_fpu_burst_8_downstream_read => nios2_fpu_burst_8_downstream_read,
      nios2_fpu_burst_8_downstream_write => nios2_fpu_burst_8_downstream_write,
      nios2_fpu_burst_8_downstream_writedata => nios2_fpu_burst_8_downstream_writedata,
      nios2_fpu_clock_0_in_endofpacket => nios2_fpu_clock_0_in_endofpacket,
      nios2_fpu_clock_0_in_readdata => nios2_fpu_clock_0_in_readdata,
      nios2_fpu_clock_0_in_waitrequest => nios2_fpu_clock_0_in_waitrequest,
      reset_n => core_clk_reset_n
    );


  --the_nios2_fpu_clock_0_out, which is an e_instance
  the_nios2_fpu_clock_0_out : nios2_fpu_clock_0_out_arbitrator
    port map(
      nios2_fpu_clock_0_out_address_to_slave => nios2_fpu_clock_0_out_address_to_slave,
      nios2_fpu_clock_0_out_endofpacket => nios2_fpu_clock_0_out_endofpacket,
      nios2_fpu_clock_0_out_readdata => nios2_fpu_clock_0_out_readdata,
      nios2_fpu_clock_0_out_reset_n => nios2_fpu_clock_0_out_reset_n,
      nios2_fpu_clock_0_out_waitrequest => nios2_fpu_clock_0_out_waitrequest,
      clk => peri_clk,
      d1_peripheral_bridge_s1_end_xfer => d1_peripheral_bridge_s1_end_xfer,
      nios2_fpu_clock_0_out_address => nios2_fpu_clock_0_out_address,
      nios2_fpu_clock_0_out_byteenable => nios2_fpu_clock_0_out_byteenable,
      nios2_fpu_clock_0_out_granted_peripheral_bridge_s1 => nios2_fpu_clock_0_out_granted_peripheral_bridge_s1,
      nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1 => nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1,
      nios2_fpu_clock_0_out_read => nios2_fpu_clock_0_out_read,
      nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1 => nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1,
      nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1_shift_register => nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1_shift_register,
      nios2_fpu_clock_0_out_requests_peripheral_bridge_s1 => nios2_fpu_clock_0_out_requests_peripheral_bridge_s1,
      nios2_fpu_clock_0_out_write => nios2_fpu_clock_0_out_write,
      nios2_fpu_clock_0_out_writedata => nios2_fpu_clock_0_out_writedata,
      peripheral_bridge_s1_endofpacket_from_sa => peripheral_bridge_s1_endofpacket_from_sa,
      peripheral_bridge_s1_readdata_from_sa => peripheral_bridge_s1_readdata_from_sa,
      peripheral_bridge_s1_waitrequest_from_sa => peripheral_bridge_s1_waitrequest_from_sa,
      reset_n => peri_clk_reset_n
    );


  --the_nios2_fpu_clock_0, which is an e_ptf_instance
  the_nios2_fpu_clock_0 : nios2_fpu_clock_0
    port map(
      master_address => nios2_fpu_clock_0_out_address,
      master_byteenable => nios2_fpu_clock_0_out_byteenable,
      master_nativeaddress => nios2_fpu_clock_0_out_nativeaddress,
      master_read => nios2_fpu_clock_0_out_read,
      master_write => nios2_fpu_clock_0_out_write,
      master_writedata => nios2_fpu_clock_0_out_writedata,
      slave_endofpacket => nios2_fpu_clock_0_in_endofpacket,
      slave_readdata => nios2_fpu_clock_0_in_readdata,
      slave_waitrequest => nios2_fpu_clock_0_in_waitrequest,
      master_clk => peri_clk,
      master_endofpacket => nios2_fpu_clock_0_out_endofpacket,
      master_readdata => nios2_fpu_clock_0_out_readdata,
      master_reset_n => nios2_fpu_clock_0_out_reset_n,
      master_waitrequest => nios2_fpu_clock_0_out_waitrequest,
      slave_address => nios2_fpu_clock_0_in_address,
      slave_byteenable => nios2_fpu_clock_0_in_byteenable,
      slave_clk => core_clk,
      slave_nativeaddress => nios2_fpu_clock_0_in_nativeaddress,
      slave_read => nios2_fpu_clock_0_in_read,
      slave_reset_n => nios2_fpu_clock_0_in_reset_n,
      slave_write => nios2_fpu_clock_0_in_write,
      slave_writedata => nios2_fpu_clock_0_in_writedata
    );


  --the_peripheral_bridge_s1, which is an e_instance
  the_peripheral_bridge_s1 : peripheral_bridge_s1_arbitrator
    port map(
      d1_peripheral_bridge_s1_end_xfer => d1_peripheral_bridge_s1_end_xfer,
      nios2_fpu_clock_0_out_granted_peripheral_bridge_s1 => nios2_fpu_clock_0_out_granted_peripheral_bridge_s1,
      nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1 => nios2_fpu_clock_0_out_qualified_request_peripheral_bridge_s1,
      nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1 => nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1,
      nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1_shift_register => nios2_fpu_clock_0_out_read_data_valid_peripheral_bridge_s1_shift_register,
      nios2_fpu_clock_0_out_requests_peripheral_bridge_s1 => nios2_fpu_clock_0_out_requests_peripheral_bridge_s1,
      peripheral_bridge_s1_address => peripheral_bridge_s1_address,
      peripheral_bridge_s1_arbiterlock => peripheral_bridge_s1_arbiterlock,
      peripheral_bridge_s1_arbiterlock2 => peripheral_bridge_s1_arbiterlock2,
      peripheral_bridge_s1_burstcount => peripheral_bridge_s1_burstcount,
      peripheral_bridge_s1_byteenable => peripheral_bridge_s1_byteenable,
      peripheral_bridge_s1_chipselect => peripheral_bridge_s1_chipselect,
      peripheral_bridge_s1_debugaccess => peripheral_bridge_s1_debugaccess,
      peripheral_bridge_s1_endofpacket_from_sa => peripheral_bridge_s1_endofpacket_from_sa,
      peripheral_bridge_s1_nativeaddress => peripheral_bridge_s1_nativeaddress,
      peripheral_bridge_s1_read => peripheral_bridge_s1_read,
      peripheral_bridge_s1_readdata_from_sa => peripheral_bridge_s1_readdata_from_sa,
      peripheral_bridge_s1_reset_n => peripheral_bridge_s1_reset_n,
      peripheral_bridge_s1_waitrequest_from_sa => peripheral_bridge_s1_waitrequest_from_sa,
      peripheral_bridge_s1_write => peripheral_bridge_s1_write,
      peripheral_bridge_s1_writedata => peripheral_bridge_s1_writedata,
      clk => peri_clk,
      nios2_fpu_clock_0_out_address_to_slave => nios2_fpu_clock_0_out_address_to_slave,
      nios2_fpu_clock_0_out_byteenable => nios2_fpu_clock_0_out_byteenable,
      nios2_fpu_clock_0_out_nativeaddress => nios2_fpu_clock_0_out_nativeaddress,
      nios2_fpu_clock_0_out_read => nios2_fpu_clock_0_out_read,
      nios2_fpu_clock_0_out_write => nios2_fpu_clock_0_out_write,
      nios2_fpu_clock_0_out_writedata => nios2_fpu_clock_0_out_writedata,
      peripheral_bridge_s1_endofpacket => peripheral_bridge_s1_endofpacket,
      peripheral_bridge_s1_readdata => peripheral_bridge_s1_readdata,
      peripheral_bridge_s1_readdatavalid => peripheral_bridge_s1_readdatavalid,
      peripheral_bridge_s1_waitrequest => peripheral_bridge_s1_waitrequest,
      reset_n => peri_clk_reset_n
    );


  --the_peripheral_bridge_m1, which is an e_instance
  the_peripheral_bridge_m1 : peripheral_bridge_m1_arbitrator
    port map(
      peripheral_bridge_m1_address_to_slave => peripheral_bridge_m1_address_to_slave,
      peripheral_bridge_m1_latency_counter => peripheral_bridge_m1_latency_counter,
      peripheral_bridge_m1_readdata => peripheral_bridge_m1_readdata,
      peripheral_bridge_m1_readdatavalid => peripheral_bridge_m1_readdatavalid,
      peripheral_bridge_m1_waitrequest => peripheral_bridge_m1_waitrequest,
      clk => peri_clk,
      d1_dipsw_s1_end_xfer => d1_dipsw_s1_end_xfer,
      d1_gpio0_s1_end_xfer => d1_gpio0_s1_end_xfer,
      d1_jtag_uart_avalon_jtag_slave_end_xfer => d1_jtag_uart_avalon_jtag_slave_end_xfer,
      d1_led_s1_end_xfer => d1_led_s1_end_xfer,
      d1_mmcdma_s1_end_xfer => d1_mmcdma_s1_end_xfer,
      d1_psw_s1_end_xfer => d1_psw_s1_end_xfer,
      d1_spu_s1_end_xfer => d1_spu_s1_end_xfer,
      d1_sysid_control_slave_end_xfer => d1_sysid_control_slave_end_xfer,
      d1_systimer_s1_end_xfer => d1_systimer_s1_end_xfer,
      d1_sysuart_s1_end_xfer => d1_sysuart_s1_end_xfer,
      d1_vga_s1_end_xfer => d1_vga_s1_end_xfer,
      dipsw_s1_readdata_from_sa => dipsw_s1_readdata_from_sa,
      gpio0_s1_readdata_from_sa => gpio0_s1_readdata_from_sa,
      jtag_uart_avalon_jtag_slave_readdata_from_sa => jtag_uart_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
      led_s1_readdata_from_sa => led_s1_readdata_from_sa,
      mmcdma_s1_readdata_from_sa => mmcdma_s1_readdata_from_sa,
      mmcdma_s1_wait_counter_eq_0 => mmcdma_s1_wait_counter_eq_0,
      peripheral_bridge_m1_address => peripheral_bridge_m1_address,
      peripheral_bridge_m1_burstcount => peripheral_bridge_m1_burstcount,
      peripheral_bridge_m1_byteenable => peripheral_bridge_m1_byteenable,
      peripheral_bridge_m1_chipselect => peripheral_bridge_m1_chipselect,
      peripheral_bridge_m1_granted_dipsw_s1 => peripheral_bridge_m1_granted_dipsw_s1,
      peripheral_bridge_m1_granted_gpio0_s1 => peripheral_bridge_m1_granted_gpio0_s1,
      peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave => peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave,
      peripheral_bridge_m1_granted_led_s1 => peripheral_bridge_m1_granted_led_s1,
      peripheral_bridge_m1_granted_mmcdma_s1 => peripheral_bridge_m1_granted_mmcdma_s1,
      peripheral_bridge_m1_granted_psw_s1 => peripheral_bridge_m1_granted_psw_s1,
      peripheral_bridge_m1_granted_spu_s1 => peripheral_bridge_m1_granted_spu_s1,
      peripheral_bridge_m1_granted_sysid_control_slave => peripheral_bridge_m1_granted_sysid_control_slave,
      peripheral_bridge_m1_granted_systimer_s1 => peripheral_bridge_m1_granted_systimer_s1,
      peripheral_bridge_m1_granted_sysuart_s1 => peripheral_bridge_m1_granted_sysuart_s1,
      peripheral_bridge_m1_granted_vga_s1 => peripheral_bridge_m1_granted_vga_s1,
      peripheral_bridge_m1_qualified_request_dipsw_s1 => peripheral_bridge_m1_qualified_request_dipsw_s1,
      peripheral_bridge_m1_qualified_request_gpio0_s1 => peripheral_bridge_m1_qualified_request_gpio0_s1,
      peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave => peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave,
      peripheral_bridge_m1_qualified_request_led_s1 => peripheral_bridge_m1_qualified_request_led_s1,
      peripheral_bridge_m1_qualified_request_mmcdma_s1 => peripheral_bridge_m1_qualified_request_mmcdma_s1,
      peripheral_bridge_m1_qualified_request_psw_s1 => peripheral_bridge_m1_qualified_request_psw_s1,
      peripheral_bridge_m1_qualified_request_spu_s1 => peripheral_bridge_m1_qualified_request_spu_s1,
      peripheral_bridge_m1_qualified_request_sysid_control_slave => peripheral_bridge_m1_qualified_request_sysid_control_slave,
      peripheral_bridge_m1_qualified_request_systimer_s1 => peripheral_bridge_m1_qualified_request_systimer_s1,
      peripheral_bridge_m1_qualified_request_sysuart_s1 => peripheral_bridge_m1_qualified_request_sysuart_s1,
      peripheral_bridge_m1_qualified_request_vga_s1 => peripheral_bridge_m1_qualified_request_vga_s1,
      peripheral_bridge_m1_read => peripheral_bridge_m1_read,
      peripheral_bridge_m1_read_data_valid_dipsw_s1 => peripheral_bridge_m1_read_data_valid_dipsw_s1,
      peripheral_bridge_m1_read_data_valid_gpio0_s1 => peripheral_bridge_m1_read_data_valid_gpio0_s1,
      peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave => peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave,
      peripheral_bridge_m1_read_data_valid_led_s1 => peripheral_bridge_m1_read_data_valid_led_s1,
      peripheral_bridge_m1_read_data_valid_mmcdma_s1 => peripheral_bridge_m1_read_data_valid_mmcdma_s1,
      peripheral_bridge_m1_read_data_valid_psw_s1 => peripheral_bridge_m1_read_data_valid_psw_s1,
      peripheral_bridge_m1_read_data_valid_spu_s1 => peripheral_bridge_m1_read_data_valid_spu_s1,
      peripheral_bridge_m1_read_data_valid_sysid_control_slave => peripheral_bridge_m1_read_data_valid_sysid_control_slave,
      peripheral_bridge_m1_read_data_valid_systimer_s1 => peripheral_bridge_m1_read_data_valid_systimer_s1,
      peripheral_bridge_m1_read_data_valid_sysuart_s1 => peripheral_bridge_m1_read_data_valid_sysuart_s1,
      peripheral_bridge_m1_read_data_valid_vga_s1 => peripheral_bridge_m1_read_data_valid_vga_s1,
      peripheral_bridge_m1_requests_dipsw_s1 => peripheral_bridge_m1_requests_dipsw_s1,
      peripheral_bridge_m1_requests_gpio0_s1 => peripheral_bridge_m1_requests_gpio0_s1,
      peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave => peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave,
      peripheral_bridge_m1_requests_led_s1 => peripheral_bridge_m1_requests_led_s1,
      peripheral_bridge_m1_requests_mmcdma_s1 => peripheral_bridge_m1_requests_mmcdma_s1,
      peripheral_bridge_m1_requests_psw_s1 => peripheral_bridge_m1_requests_psw_s1,
      peripheral_bridge_m1_requests_spu_s1 => peripheral_bridge_m1_requests_spu_s1,
      peripheral_bridge_m1_requests_sysid_control_slave => peripheral_bridge_m1_requests_sysid_control_slave,
      peripheral_bridge_m1_requests_systimer_s1 => peripheral_bridge_m1_requests_systimer_s1,
      peripheral_bridge_m1_requests_sysuart_s1 => peripheral_bridge_m1_requests_sysuart_s1,
      peripheral_bridge_m1_requests_vga_s1 => peripheral_bridge_m1_requests_vga_s1,
      peripheral_bridge_m1_write => peripheral_bridge_m1_write,
      peripheral_bridge_m1_writedata => peripheral_bridge_m1_writedata,
      psw_s1_readdata_from_sa => psw_s1_readdata_from_sa,
      reset_n => peri_clk_reset_n,
      spu_s1_readdata_from_sa => spu_s1_readdata_from_sa,
      spu_s1_waitrequest_from_sa => spu_s1_waitrequest_from_sa,
      sysid_control_slave_readdata_from_sa => sysid_control_slave_readdata_from_sa,
      systimer_s1_readdata_from_sa => systimer_s1_readdata_from_sa,
      sysuart_s1_readdata_from_sa => sysuart_s1_readdata_from_sa,
      vga_s1_readdata_from_sa => vga_s1_readdata_from_sa
    );


  --the_peripheral_bridge, which is an e_ptf_instance
  the_peripheral_bridge : peripheral_bridge
    port map(
      m1_address => peripheral_bridge_m1_address,
      m1_burstcount => peripheral_bridge_m1_burstcount,
      m1_byteenable => peripheral_bridge_m1_byteenable,
      m1_chipselect => peripheral_bridge_m1_chipselect,
      m1_debugaccess => peripheral_bridge_m1_debugaccess,
      m1_read => peripheral_bridge_m1_read,
      m1_write => peripheral_bridge_m1_write,
      m1_writedata => peripheral_bridge_m1_writedata,
      s1_endofpacket => peripheral_bridge_s1_endofpacket,
      s1_readdata => peripheral_bridge_s1_readdata,
      s1_readdatavalid => peripheral_bridge_s1_readdatavalid,
      s1_waitrequest => peripheral_bridge_s1_waitrequest,
      clk => peri_clk,
      m1_endofpacket => peripheral_bridge_m1_endofpacket,
      m1_readdata => peripheral_bridge_m1_readdata,
      m1_readdatavalid => peripheral_bridge_m1_readdatavalid,
      m1_waitrequest => peripheral_bridge_m1_waitrequest,
      reset_n => peripheral_bridge_s1_reset_n,
      s1_address => peripheral_bridge_s1_address,
      s1_arbiterlock => peripheral_bridge_s1_arbiterlock,
      s1_arbiterlock2 => peripheral_bridge_s1_arbiterlock2,
      s1_burstcount => peripheral_bridge_s1_burstcount,
      s1_byteenable => peripheral_bridge_s1_byteenable,
      s1_chipselect => peripheral_bridge_s1_chipselect,
      s1_debugaccess => peripheral_bridge_s1_debugaccess,
      s1_nativeaddress => peripheral_bridge_s1_nativeaddress,
      s1_read => peripheral_bridge_s1_read,
      s1_write => peripheral_bridge_s1_write,
      s1_writedata => peripheral_bridge_s1_writedata
    );


  --the_psw_s1, which is an e_instance
  the_psw_s1 : psw_s1_arbitrator
    port map(
      d1_psw_s1_end_xfer => d1_psw_s1_end_xfer,
      peripheral_bridge_m1_granted_psw_s1 => peripheral_bridge_m1_granted_psw_s1,
      peripheral_bridge_m1_qualified_request_psw_s1 => peripheral_bridge_m1_qualified_request_psw_s1,
      peripheral_bridge_m1_read_data_valid_psw_s1 => peripheral_bridge_m1_read_data_valid_psw_s1,
      peripheral_bridge_m1_requests_psw_s1 => peripheral_bridge_m1_requests_psw_s1,
      psw_s1_address => psw_s1_address,
      psw_s1_chipselect => psw_s1_chipselect,
      psw_s1_irq_from_sa => psw_s1_irq_from_sa,
      psw_s1_readdata_from_sa => psw_s1_readdata_from_sa,
      psw_s1_reset_n => psw_s1_reset_n,
      psw_s1_write_n => psw_s1_write_n,
      psw_s1_writedata => psw_s1_writedata,
      clk => peri_clk,
      peripheral_bridge_m1_address_to_slave => peripheral_bridge_m1_address_to_slave,
      peripheral_bridge_m1_burstcount => peripheral_bridge_m1_burstcount,
      peripheral_bridge_m1_chipselect => peripheral_bridge_m1_chipselect,
      peripheral_bridge_m1_latency_counter => peripheral_bridge_m1_latency_counter,
      peripheral_bridge_m1_read => peripheral_bridge_m1_read,
      peripheral_bridge_m1_write => peripheral_bridge_m1_write,
      peripheral_bridge_m1_writedata => peripheral_bridge_m1_writedata,
      psw_s1_irq => psw_s1_irq,
      psw_s1_readdata => psw_s1_readdata,
      reset_n => peri_clk_reset_n
    );


  --the_psw, which is an e_ptf_instance
  the_psw : psw
    port map(
      irq => psw_s1_irq,
      readdata => psw_s1_readdata,
      address => psw_s1_address,
      chipselect => psw_s1_chipselect,
      clk => peri_clk,
      in_port => in_port_to_the_psw,
      reset_n => psw_s1_reset_n,
      write_n => psw_s1_write_n,
      writedata => psw_s1_writedata
    );


  --the_sdram_s1, which is an e_instance
  the_sdram_s1 : sdram_s1_arbitrator
    port map(
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      nios2_fpu_burst_0_downstream_granted_sdram_s1 => nios2_fpu_burst_0_downstream_granted_sdram_s1,
      nios2_fpu_burst_0_downstream_qualified_request_sdram_s1 => nios2_fpu_burst_0_downstream_qualified_request_sdram_s1,
      nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1 => nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1,
      nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1_shift_register => nios2_fpu_burst_0_downstream_read_data_valid_sdram_s1_shift_register,
      nios2_fpu_burst_0_downstream_requests_sdram_s1 => nios2_fpu_burst_0_downstream_requests_sdram_s1,
      nios2_fpu_burst_1_downstream_granted_sdram_s1 => nios2_fpu_burst_1_downstream_granted_sdram_s1,
      nios2_fpu_burst_1_downstream_qualified_request_sdram_s1 => nios2_fpu_burst_1_downstream_qualified_request_sdram_s1,
      nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1 => nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1,
      nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1_shift_register => nios2_fpu_burst_1_downstream_read_data_valid_sdram_s1_shift_register,
      nios2_fpu_burst_1_downstream_requests_sdram_s1 => nios2_fpu_burst_1_downstream_requests_sdram_s1,
      nios2_fpu_burst_2_downstream_granted_sdram_s1 => nios2_fpu_burst_2_downstream_granted_sdram_s1,
      nios2_fpu_burst_2_downstream_qualified_request_sdram_s1 => nios2_fpu_burst_2_downstream_qualified_request_sdram_s1,
      nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1 => nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1,
      nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1_shift_register => nios2_fpu_burst_2_downstream_read_data_valid_sdram_s1_shift_register,
      nios2_fpu_burst_2_downstream_requests_sdram_s1 => nios2_fpu_burst_2_downstream_requests_sdram_s1,
      nios2_fpu_burst_3_downstream_granted_sdram_s1 => nios2_fpu_burst_3_downstream_granted_sdram_s1,
      nios2_fpu_burst_3_downstream_qualified_request_sdram_s1 => nios2_fpu_burst_3_downstream_qualified_request_sdram_s1,
      nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1 => nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1,
      nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1_shift_register => nios2_fpu_burst_3_downstream_read_data_valid_sdram_s1_shift_register,
      nios2_fpu_burst_3_downstream_requests_sdram_s1 => nios2_fpu_burst_3_downstream_requests_sdram_s1,
      sdram_s1_address => sdram_s1_address,
      sdram_s1_byteenable_n => sdram_s1_byteenable_n,
      sdram_s1_chipselect => sdram_s1_chipselect,
      sdram_s1_read_n => sdram_s1_read_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_reset_n => sdram_s1_reset_n,
      sdram_s1_waitrequest_from_sa => sdram_s1_waitrequest_from_sa,
      sdram_s1_write_n => sdram_s1_write_n,
      sdram_s1_writedata => sdram_s1_writedata,
      clk => core_clk,
      nios2_fpu_burst_0_downstream_address_to_slave => nios2_fpu_burst_0_downstream_address_to_slave,
      nios2_fpu_burst_0_downstream_arbitrationshare => nios2_fpu_burst_0_downstream_arbitrationshare,
      nios2_fpu_burst_0_downstream_burstcount => nios2_fpu_burst_0_downstream_burstcount,
      nios2_fpu_burst_0_downstream_byteenable => nios2_fpu_burst_0_downstream_byteenable,
      nios2_fpu_burst_0_downstream_latency_counter => nios2_fpu_burst_0_downstream_latency_counter,
      nios2_fpu_burst_0_downstream_read => nios2_fpu_burst_0_downstream_read,
      nios2_fpu_burst_0_downstream_write => nios2_fpu_burst_0_downstream_write,
      nios2_fpu_burst_0_downstream_writedata => nios2_fpu_burst_0_downstream_writedata,
      nios2_fpu_burst_1_downstream_address_to_slave => nios2_fpu_burst_1_downstream_address_to_slave,
      nios2_fpu_burst_1_downstream_arbitrationshare => nios2_fpu_burst_1_downstream_arbitrationshare,
      nios2_fpu_burst_1_downstream_burstcount => nios2_fpu_burst_1_downstream_burstcount,
      nios2_fpu_burst_1_downstream_byteenable => nios2_fpu_burst_1_downstream_byteenable,
      nios2_fpu_burst_1_downstream_latency_counter => nios2_fpu_burst_1_downstream_latency_counter,
      nios2_fpu_burst_1_downstream_read => nios2_fpu_burst_1_downstream_read,
      nios2_fpu_burst_1_downstream_write => nios2_fpu_burst_1_downstream_write,
      nios2_fpu_burst_1_downstream_writedata => nios2_fpu_burst_1_downstream_writedata,
      nios2_fpu_burst_2_downstream_address_to_slave => nios2_fpu_burst_2_downstream_address_to_slave,
      nios2_fpu_burst_2_downstream_arbitrationshare => nios2_fpu_burst_2_downstream_arbitrationshare,
      nios2_fpu_burst_2_downstream_burstcount => nios2_fpu_burst_2_downstream_burstcount,
      nios2_fpu_burst_2_downstream_byteenable => nios2_fpu_burst_2_downstream_byteenable,
      nios2_fpu_burst_2_downstream_latency_counter => nios2_fpu_burst_2_downstream_latency_counter,
      nios2_fpu_burst_2_downstream_read => nios2_fpu_burst_2_downstream_read,
      nios2_fpu_burst_2_downstream_write => nios2_fpu_burst_2_downstream_write,
      nios2_fpu_burst_2_downstream_writedata => nios2_fpu_burst_2_downstream_writedata,
      nios2_fpu_burst_3_downstream_address_to_slave => nios2_fpu_burst_3_downstream_address_to_slave,
      nios2_fpu_burst_3_downstream_arbitrationshare => nios2_fpu_burst_3_downstream_arbitrationshare,
      nios2_fpu_burst_3_downstream_burstcount => nios2_fpu_burst_3_downstream_burstcount,
      nios2_fpu_burst_3_downstream_byteenable => nios2_fpu_burst_3_downstream_byteenable,
      nios2_fpu_burst_3_downstream_latency_counter => nios2_fpu_burst_3_downstream_latency_counter,
      nios2_fpu_burst_3_downstream_read => nios2_fpu_burst_3_downstream_read,
      nios2_fpu_burst_3_downstream_write => nios2_fpu_burst_3_downstream_write,
      nios2_fpu_burst_3_downstream_writedata => nios2_fpu_burst_3_downstream_writedata,
      reset_n => core_clk_reset_n,
      sdram_s1_readdata => sdram_s1_readdata,
      sdram_s1_readdatavalid => sdram_s1_readdatavalid,
      sdram_s1_waitrequest => sdram_s1_waitrequest
    );


  --the_sdram, which is an e_ptf_instance
  the_sdram : sdram
    port map(
      za_data => sdram_s1_readdata,
      za_valid => sdram_s1_readdatavalid,
      za_waitrequest => sdram_s1_waitrequest,
      zs_addr => internal_zs_addr_from_the_sdram,
      zs_ba => internal_zs_ba_from_the_sdram,
      zs_cas_n => internal_zs_cas_n_from_the_sdram,
      zs_cke => internal_zs_cke_from_the_sdram,
      zs_cs_n => internal_zs_cs_n_from_the_sdram,
      zs_dq => zs_dq_to_and_from_the_sdram,
      zs_dqm => internal_zs_dqm_from_the_sdram,
      zs_ras_n => internal_zs_ras_n_from_the_sdram,
      zs_we_n => internal_zs_we_n_from_the_sdram,
      az_addr => sdram_s1_address,
      az_be_n => sdram_s1_byteenable_n,
      az_cs => sdram_s1_chipselect,
      az_data => sdram_s1_writedata,
      az_rd_n => sdram_s1_read_n,
      az_wr_n => sdram_s1_write_n,
      clk => core_clk,
      reset_n => sdram_s1_reset_n
    );


  --the_spu_s1, which is an e_instance
  the_spu_s1 : spu_s1_arbitrator
    port map(
      d1_spu_s1_end_xfer => d1_spu_s1_end_xfer,
      peripheral_bridge_m1_granted_spu_s1 => peripheral_bridge_m1_granted_spu_s1,
      peripheral_bridge_m1_qualified_request_spu_s1 => peripheral_bridge_m1_qualified_request_spu_s1,
      peripheral_bridge_m1_read_data_valid_spu_s1 => peripheral_bridge_m1_read_data_valid_spu_s1,
      peripheral_bridge_m1_requests_spu_s1 => peripheral_bridge_m1_requests_spu_s1,
      spu_s1_address => spu_s1_address,
      spu_s1_byteenable => spu_s1_byteenable,
      spu_s1_chipselect => spu_s1_chipselect,
      spu_s1_irq_from_sa => spu_s1_irq_from_sa,
      spu_s1_read => spu_s1_read,
      spu_s1_readdata_from_sa => spu_s1_readdata_from_sa,
      spu_s1_reset => spu_s1_reset,
      spu_s1_waitrequest_from_sa => spu_s1_waitrequest_from_sa,
      spu_s1_write => spu_s1_write,
      spu_s1_writedata => spu_s1_writedata,
      clk => peri_clk,
      peripheral_bridge_m1_address_to_slave => peripheral_bridge_m1_address_to_slave,
      peripheral_bridge_m1_burstcount => peripheral_bridge_m1_burstcount,
      peripheral_bridge_m1_byteenable => peripheral_bridge_m1_byteenable,
      peripheral_bridge_m1_chipselect => peripheral_bridge_m1_chipselect,
      peripheral_bridge_m1_latency_counter => peripheral_bridge_m1_latency_counter,
      peripheral_bridge_m1_read => peripheral_bridge_m1_read,
      peripheral_bridge_m1_write => peripheral_bridge_m1_write,
      peripheral_bridge_m1_writedata => peripheral_bridge_m1_writedata,
      reset_n => peri_clk_reset_n,
      spu_s1_irq => spu_s1_irq,
      spu_s1_readdata => spu_s1_readdata,
      spu_s1_waitrequest => spu_s1_waitrequest
    );


  --the_spu_m1, which is an e_instance
  the_spu_m1 : spu_m1_arbitrator
    port map(
      spu_m1_address_to_slave => spu_m1_address_to_slave,
      spu_m1_latency_counter => spu_m1_latency_counter,
      spu_m1_readdata => spu_m1_readdata,
      spu_m1_readdatavalid => spu_m1_readdatavalid,
      spu_m1_waitrequest => spu_m1_waitrequest,
      clk => core_clk,
      d1_nios2_fpu_burst_3_upstream_end_xfer => d1_nios2_fpu_burst_3_upstream_end_xfer,
      nios2_fpu_burst_3_upstream_readdata_from_sa => nios2_fpu_burst_3_upstream_readdata_from_sa,
      nios2_fpu_burst_3_upstream_waitrequest_from_sa => nios2_fpu_burst_3_upstream_waitrequest_from_sa,
      reset_n => core_clk_reset_n,
      spu_m1_address => spu_m1_address,
      spu_m1_burstcount => spu_m1_burstcount,
      spu_m1_granted_nios2_fpu_burst_3_upstream => spu_m1_granted_nios2_fpu_burst_3_upstream,
      spu_m1_qualified_request_nios2_fpu_burst_3_upstream => spu_m1_qualified_request_nios2_fpu_burst_3_upstream,
      spu_m1_read => spu_m1_read,
      spu_m1_read_data_valid_nios2_fpu_burst_3_upstream => spu_m1_read_data_valid_nios2_fpu_burst_3_upstream,
      spu_m1_read_data_valid_nios2_fpu_burst_3_upstream_shift_register => spu_m1_read_data_valid_nios2_fpu_burst_3_upstream_shift_register,
      spu_m1_requests_nios2_fpu_burst_3_upstream => spu_m1_requests_nios2_fpu_burst_3_upstream
    );


  --the_spu, which is an e_ptf_instance
  the_spu : spu
    port map(
      AUD_L => internal_AUD_L_from_the_spu,
      AUD_R => internal_AUD_R_from_the_spu,
      DAC_BCLK => internal_DAC_BCLK_from_the_spu,
      DAC_DATA => internal_DAC_DATA_from_the_spu,
      DAC_LRCK => internal_DAC_LRCK_from_the_spu,
      SPDIF => internal_SPDIF_from_the_spu,
      avm_m1_address => spu_m1_address,
      avm_m1_burstcount => spu_m1_burstcount,
      avm_m1_read => spu_m1_read,
      avs_s1_irq => spu_s1_irq,
      avs_s1_readdata => spu_s1_readdata,
      avs_s1_waitrequest => spu_s1_waitrequest,
      avm_m1_readdata => spu_m1_readdata,
      avm_m1_readdatavalid => spu_m1_readdatavalid,
      avm_m1_waitrequest => spu_m1_waitrequest,
      avs_s1_address => spu_s1_address,
      avs_s1_byteenable => spu_s1_byteenable,
      avs_s1_chipselect => spu_s1_chipselect,
      avs_s1_read => spu_s1_read,
      avs_s1_write => spu_s1_write,
      avs_s1_writedata => spu_s1_writedata,
      clk_128fs => clk_128fs_to_the_spu,
      csi_global_clock => peri_clk,
      csi_global_reset => spu_s1_reset,
      csi_m1_clock => core_clk
    );


  --the_sysid_control_slave, which is an e_instance
  the_sysid_control_slave : sysid_control_slave_arbitrator
    port map(
      d1_sysid_control_slave_end_xfer => d1_sysid_control_slave_end_xfer,
      peripheral_bridge_m1_granted_sysid_control_slave => peripheral_bridge_m1_granted_sysid_control_slave,
      peripheral_bridge_m1_qualified_request_sysid_control_slave => peripheral_bridge_m1_qualified_request_sysid_control_slave,
      peripheral_bridge_m1_read_data_valid_sysid_control_slave => peripheral_bridge_m1_read_data_valid_sysid_control_slave,
      peripheral_bridge_m1_requests_sysid_control_slave => peripheral_bridge_m1_requests_sysid_control_slave,
      sysid_control_slave_address => sysid_control_slave_address,
      sysid_control_slave_readdata_from_sa => sysid_control_slave_readdata_from_sa,
      sysid_control_slave_reset_n => sysid_control_slave_reset_n,
      clk => peri_clk,
      peripheral_bridge_m1_address_to_slave => peripheral_bridge_m1_address_to_slave,
      peripheral_bridge_m1_burstcount => peripheral_bridge_m1_burstcount,
      peripheral_bridge_m1_chipselect => peripheral_bridge_m1_chipselect,
      peripheral_bridge_m1_latency_counter => peripheral_bridge_m1_latency_counter,
      peripheral_bridge_m1_read => peripheral_bridge_m1_read,
      peripheral_bridge_m1_write => peripheral_bridge_m1_write,
      reset_n => peri_clk_reset_n,
      sysid_control_slave_readdata => sysid_control_slave_readdata
    );


  --the_sysid, which is an e_ptf_instance
  the_sysid : sysid
    port map(
      readdata => sysid_control_slave_readdata,
      address => sysid_control_slave_address,
      clock => sysid_control_slave_clock,
      reset_n => sysid_control_slave_reset_n
    );


  --the_systimer_s1, which is an e_instance
  the_systimer_s1 : systimer_s1_arbitrator
    port map(
      d1_systimer_s1_end_xfer => d1_systimer_s1_end_xfer,
      peripheral_bridge_m1_granted_systimer_s1 => peripheral_bridge_m1_granted_systimer_s1,
      peripheral_bridge_m1_qualified_request_systimer_s1 => peripheral_bridge_m1_qualified_request_systimer_s1,
      peripheral_bridge_m1_read_data_valid_systimer_s1 => peripheral_bridge_m1_read_data_valid_systimer_s1,
      peripheral_bridge_m1_requests_systimer_s1 => peripheral_bridge_m1_requests_systimer_s1,
      systimer_s1_address => systimer_s1_address,
      systimer_s1_chipselect => systimer_s1_chipselect,
      systimer_s1_irq_from_sa => systimer_s1_irq_from_sa,
      systimer_s1_readdata_from_sa => systimer_s1_readdata_from_sa,
      systimer_s1_reset_n => systimer_s1_reset_n,
      systimer_s1_write_n => systimer_s1_write_n,
      systimer_s1_writedata => systimer_s1_writedata,
      clk => peri_clk,
      peripheral_bridge_m1_address_to_slave => peripheral_bridge_m1_address_to_slave,
      peripheral_bridge_m1_burstcount => peripheral_bridge_m1_burstcount,
      peripheral_bridge_m1_chipselect => peripheral_bridge_m1_chipselect,
      peripheral_bridge_m1_latency_counter => peripheral_bridge_m1_latency_counter,
      peripheral_bridge_m1_read => peripheral_bridge_m1_read,
      peripheral_bridge_m1_write => peripheral_bridge_m1_write,
      peripheral_bridge_m1_writedata => peripheral_bridge_m1_writedata,
      reset_n => peri_clk_reset_n,
      systimer_s1_irq => systimer_s1_irq,
      systimer_s1_readdata => systimer_s1_readdata
    );


  --the_systimer, which is an e_ptf_instance
  the_systimer : systimer
    port map(
      irq => systimer_s1_irq,
      readdata => systimer_s1_readdata,
      address => systimer_s1_address,
      chipselect => systimer_s1_chipselect,
      clk => peri_clk,
      reset_n => systimer_s1_reset_n,
      write_n => systimer_s1_write_n,
      writedata => systimer_s1_writedata
    );


  --the_sysuart_s1, which is an e_instance
  the_sysuart_s1 : sysuart_s1_arbitrator
    port map(
      d1_sysuart_s1_end_xfer => d1_sysuart_s1_end_xfer,
      peripheral_bridge_m1_granted_sysuart_s1 => peripheral_bridge_m1_granted_sysuart_s1,
      peripheral_bridge_m1_qualified_request_sysuart_s1 => peripheral_bridge_m1_qualified_request_sysuart_s1,
      peripheral_bridge_m1_read_data_valid_sysuart_s1 => peripheral_bridge_m1_read_data_valid_sysuart_s1,
      peripheral_bridge_m1_requests_sysuart_s1 => peripheral_bridge_m1_requests_sysuart_s1,
      sysuart_s1_address => sysuart_s1_address,
      sysuart_s1_begintransfer => sysuart_s1_begintransfer,
      sysuart_s1_chipselect => sysuart_s1_chipselect,
      sysuart_s1_dataavailable_from_sa => sysuart_s1_dataavailable_from_sa,
      sysuart_s1_irq_from_sa => sysuart_s1_irq_from_sa,
      sysuart_s1_read_n => sysuart_s1_read_n,
      sysuart_s1_readdata_from_sa => sysuart_s1_readdata_from_sa,
      sysuart_s1_readyfordata_from_sa => sysuart_s1_readyfordata_from_sa,
      sysuart_s1_reset_n => sysuart_s1_reset_n,
      sysuart_s1_write_n => sysuart_s1_write_n,
      sysuart_s1_writedata => sysuart_s1_writedata,
      clk => peri_clk,
      peripheral_bridge_m1_address_to_slave => peripheral_bridge_m1_address_to_slave,
      peripheral_bridge_m1_burstcount => peripheral_bridge_m1_burstcount,
      peripheral_bridge_m1_chipselect => peripheral_bridge_m1_chipselect,
      peripheral_bridge_m1_latency_counter => peripheral_bridge_m1_latency_counter,
      peripheral_bridge_m1_read => peripheral_bridge_m1_read,
      peripheral_bridge_m1_write => peripheral_bridge_m1_write,
      peripheral_bridge_m1_writedata => peripheral_bridge_m1_writedata,
      reset_n => peri_clk_reset_n,
      sysuart_s1_dataavailable => sysuart_s1_dataavailable,
      sysuart_s1_irq => sysuart_s1_irq,
      sysuart_s1_readdata => sysuart_s1_readdata,
      sysuart_s1_readyfordata => sysuart_s1_readyfordata
    );


  --the_sysuart, which is an e_ptf_instance
  the_sysuart : sysuart
    port map(
      dataavailable => sysuart_s1_dataavailable,
      irq => sysuart_s1_irq,
      readdata => sysuart_s1_readdata,
      readyfordata => sysuart_s1_readyfordata,
      txd => internal_txd_from_the_sysuart,
      address => sysuart_s1_address,
      begintransfer => sysuart_s1_begintransfer,
      chipselect => sysuart_s1_chipselect,
      clk => peri_clk,
      read_n => sysuart_s1_read_n,
      reset_n => sysuart_s1_reset_n,
      rxd => rxd_to_the_sysuart,
      write_n => sysuart_s1_write_n,
      writedata => sysuart_s1_writedata
    );


  --the_vga_s1, which is an e_instance
  the_vga_s1 : vga_s1_arbitrator
    port map(
      d1_vga_s1_end_xfer => d1_vga_s1_end_xfer,
      peripheral_bridge_m1_granted_vga_s1 => peripheral_bridge_m1_granted_vga_s1,
      peripheral_bridge_m1_qualified_request_vga_s1 => peripheral_bridge_m1_qualified_request_vga_s1,
      peripheral_bridge_m1_read_data_valid_vga_s1 => peripheral_bridge_m1_read_data_valid_vga_s1,
      peripheral_bridge_m1_requests_vga_s1 => peripheral_bridge_m1_requests_vga_s1,
      vga_s1_address => vga_s1_address,
      vga_s1_irq_from_sa => vga_s1_irq_from_sa,
      vga_s1_read => vga_s1_read,
      vga_s1_readdata_from_sa => vga_s1_readdata_from_sa,
      vga_s1_write => vga_s1_write,
      vga_s1_writedata => vga_s1_writedata,
      clk => peri_clk,
      peripheral_bridge_m1_address_to_slave => peripheral_bridge_m1_address_to_slave,
      peripheral_bridge_m1_burstcount => peripheral_bridge_m1_burstcount,
      peripheral_bridge_m1_chipselect => peripheral_bridge_m1_chipselect,
      peripheral_bridge_m1_latency_counter => peripheral_bridge_m1_latency_counter,
      peripheral_bridge_m1_read => peripheral_bridge_m1_read,
      peripheral_bridge_m1_write => peripheral_bridge_m1_write,
      peripheral_bridge_m1_writedata => peripheral_bridge_m1_writedata,
      reset_n => peri_clk_reset_n,
      vga_s1_irq => vga_s1_irq,
      vga_s1_readdata => vga_s1_readdata
    );


  --the_vga_m1, which is an e_instance
  the_vga_m1 : vga_m1_arbitrator
    port map(
      vga_m1_address_to_slave => vga_m1_address_to_slave,
      vga_m1_dbs_address => vga_m1_dbs_address,
      vga_m1_latency_counter => vga_m1_latency_counter,
      vga_m1_readdata => vga_m1_readdata,
      vga_m1_readdatavalid => vga_m1_readdatavalid,
      vga_m1_reset => vga_m1_reset,
      vga_m1_waitrequest => vga_m1_waitrequest,
      clk => core_clk,
      d1_nios2_fpu_burst_0_upstream_end_xfer => d1_nios2_fpu_burst_0_upstream_end_xfer,
      nios2_fpu_burst_0_upstream_readdata_from_sa => nios2_fpu_burst_0_upstream_readdata_from_sa,
      nios2_fpu_burst_0_upstream_waitrequest_from_sa => nios2_fpu_burst_0_upstream_waitrequest_from_sa,
      reset_n => core_clk_reset_n,
      vga_m1_address => vga_m1_address,
      vga_m1_burstcount => vga_m1_burstcount,
      vga_m1_granted_nios2_fpu_burst_0_upstream => vga_m1_granted_nios2_fpu_burst_0_upstream,
      vga_m1_qualified_request_nios2_fpu_burst_0_upstream => vga_m1_qualified_request_nios2_fpu_burst_0_upstream,
      vga_m1_read => vga_m1_read,
      vga_m1_read_data_valid_nios2_fpu_burst_0_upstream => vga_m1_read_data_valid_nios2_fpu_burst_0_upstream,
      vga_m1_read_data_valid_nios2_fpu_burst_0_upstream_shift_register => vga_m1_read_data_valid_nios2_fpu_burst_0_upstream_shift_register,
      vga_m1_requests_nios2_fpu_burst_0_upstream => vga_m1_requests_nios2_fpu_burst_0_upstream
    );


  --the_vga, which is an e_ptf_instance
  the_vga : vga
    port map(
      avm_m1_address => vga_m1_address,
      avm_m1_burstcount => vga_m1_burstcount,
      avm_m1_read => vga_m1_read,
      avs_s1_readdata => vga_s1_readdata,
      irq_s1 => vga_s1_irq,
      video_bout => internal_video_bout_from_the_vga,
      video_enable => internal_video_enable_from_the_vga,
      video_gout => internal_video_gout_from_the_vga,
      video_hsync_n => internal_video_hsync_n_from_the_vga,
      video_rout => internal_video_rout_from_the_vga,
      video_vsync_n => internal_video_vsync_n_from_the_vga,
      avm_m1_readdata => vga_m1_readdata,
      avm_m1_readdatavalid => vga_m1_readdatavalid,
      avm_m1_waitrequest => vga_m1_waitrequest,
      avs_s1_address => vga_s1_address,
      avs_s1_read => vga_s1_read,
      avs_s1_write => vga_s1_write,
      avs_s1_writedata => vga_s1_writedata,
      csi_m1_clk => core_clk,
      csi_m1_reset => vga_m1_reset,
      csi_s1_clk => peri_clk,
      video_clk => video_clk_to_the_vga
    );


  --reset is asserted asynchronously and deasserted synchronously
  nios2_fpu_reset_peri_clk_domain_synch : nios2_fpu_reset_peri_clk_domain_synch_module
    port map(
      data_out => peri_clk_reset_n,
      clk => peri_clk,
      data_in => module_input69,
      reset_n => reset_n_sources
    );

  module_input69 <= std_logic'('1');

  --reset sources mux, which is an e_mux
  reset_n_sources <= Vector_To_Std_Logic(NOT ((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT reset_n))) OR std_logic_vector'("00000000000000000000000000000000")) OR std_logic_vector'("00000000000000000000000000000000")) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_jtag_debug_module_resetrequest_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(nios2_fast_fpu_jtag_debug_module_resetrequest_from_sa))))));
  --reset is asserted asynchronously and deasserted synchronously
  nios2_fpu_reset_core_clk_domain_synch : nios2_fpu_reset_core_clk_domain_synch_module
    port map(
      data_out => core_clk_reset_n,
      clk => core_clk,
      data_in => module_input70,
      reset_n => reset_n_sources
    );

  module_input70 <= std_logic'('1');

  --nios2_fpu_burst_0_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  nios2_fpu_burst_0_upstream_writedata <= std_logic_vector'("0000000000000000");
  --nios2_fpu_burst_1_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  nios2_fpu_burst_1_upstream_writedata <= std_logic_vector'("0000000000000000");
  --nios2_fpu_burst_3_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  nios2_fpu_burst_3_upstream_writedata <= std_logic_vector'("0000000000000000");
  --nios2_fpu_burst_4_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  nios2_fpu_burst_4_upstream_writedata <= std_logic_vector'("00000000000000000000000000000000");
  --nios2_fpu_burst_7_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  nios2_fpu_burst_7_upstream_writedata <= std_logic_vector'("00000000000000000000000000000000");
  --peripheral_bridge_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  peripheral_bridge_m1_endofpacket <= std_logic'('0');
  --sysid_control_slave_clock of type clock does not connect to anything so wire it to default (0)
  sysid_control_slave_clock <= std_logic'('0');
  --vhdl renameroo for output signals
  AUD_L_from_the_spu <= internal_AUD_L_from_the_spu;
  --vhdl renameroo for output signals
  AUD_R_from_the_spu <= internal_AUD_R_from_the_spu;
  --vhdl renameroo for output signals
  DAC_BCLK_from_the_spu <= internal_DAC_BCLK_from_the_spu;
  --vhdl renameroo for output signals
  DAC_DATA_from_the_spu <= internal_DAC_DATA_from_the_spu;
  --vhdl renameroo for output signals
  DAC_LRCK_from_the_spu <= internal_DAC_LRCK_from_the_spu;
  --vhdl renameroo for output signals
  MMC_SCK_from_the_mmcdma <= internal_MMC_SCK_from_the_mmcdma;
  --vhdl renameroo for output signals
  MMC_SDO_from_the_mmcdma <= internal_MMC_SDO_from_the_mmcdma;
  --vhdl renameroo for output signals
  MMC_nCS_from_the_mmcdma <= internal_MMC_nCS_from_the_mmcdma;
  --vhdl renameroo for output signals
  SPDIF_from_the_spu <= internal_SPDIF_from_the_spu;
  --vhdl renameroo for output signals
  out_port_from_the_led <= internal_out_port_from_the_led;
  --vhdl renameroo for output signals
  txd_from_the_sysuart <= internal_txd_from_the_sysuart;
  --vhdl renameroo for output signals
  video_bout_from_the_vga <= internal_video_bout_from_the_vga;
  --vhdl renameroo for output signals
  video_enable_from_the_vga <= internal_video_enable_from_the_vga;
  --vhdl renameroo for output signals
  video_gout_from_the_vga <= internal_video_gout_from_the_vga;
  --vhdl renameroo for output signals
  video_hsync_n_from_the_vga <= internal_video_hsync_n_from_the_vga;
  --vhdl renameroo for output signals
  video_rout_from_the_vga <= internal_video_rout_from_the_vga;
  --vhdl renameroo for output signals
  video_vsync_n_from_the_vga <= internal_video_vsync_n_from_the_vga;
  --vhdl renameroo for output signals
  zs_addr_from_the_sdram <= internal_zs_addr_from_the_sdram;
  --vhdl renameroo for output signals
  zs_ba_from_the_sdram <= internal_zs_ba_from_the_sdram;
  --vhdl renameroo for output signals
  zs_cas_n_from_the_sdram <= internal_zs_cas_n_from_the_sdram;
  --vhdl renameroo for output signals
  zs_cke_from_the_sdram <= internal_zs_cke_from_the_sdram;
  --vhdl renameroo for output signals
  zs_cs_n_from_the_sdram <= internal_zs_cs_n_from_the_sdram;
  --vhdl renameroo for output signals
  zs_dqm_from_the_sdram <= internal_zs_dqm_from_the_sdram;
  --vhdl renameroo for output signals
  zs_ras_n_from_the_sdram <= internal_zs_ras_n_from_the_sdram;
  --vhdl renameroo for output signals
  zs_we_n_from_the_sdram <= internal_zs_we_n_from_the_sdram;

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library altera_mf;
use altera_mf.altera_mf_components.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;



-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your libraries here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>

entity test_bench is 
end entity test_bench;


architecture europa of test_bench is
component nios2_fpu is 
           port (
                 -- 1) global signals:
                    signal core_clk : IN STD_LOGIC;
                    signal peri_clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- the_dipsw
                    signal in_port_to_the_dipsw : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- the_gpio0
                    signal bidir_port_to_and_from_the_gpio0 : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- the_led
                    signal out_port_from_the_led : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_mmcdma
                    signal MMC_CD_to_the_mmcdma : IN STD_LOGIC;
                    signal MMC_SCK_from_the_mmcdma : OUT STD_LOGIC;
                    signal MMC_SDI_to_the_mmcdma : IN STD_LOGIC;
                    signal MMC_SDO_from_the_mmcdma : OUT STD_LOGIC;
                    signal MMC_WP_to_the_mmcdma : IN STD_LOGIC;
                    signal MMC_nCS_from_the_mmcdma : OUT STD_LOGIC;

                 -- the_psw
                    signal in_port_to_the_psw : IN STD_LOGIC_VECTOR (1 DOWNTO 0);

                 -- the_sdram
                    signal zs_addr_from_the_sdram : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal zs_ba_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_cas_n_from_the_sdram : OUT STD_LOGIC;
                    signal zs_cke_from_the_sdram : OUT STD_LOGIC;
                    signal zs_cs_n_from_the_sdram : OUT STD_LOGIC;
                    signal zs_dq_to_and_from_the_sdram : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal zs_dqm_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_ras_n_from_the_sdram : OUT STD_LOGIC;
                    signal zs_we_n_from_the_sdram : OUT STD_LOGIC;

                 -- the_spu
                    signal AUD_L_from_the_spu : OUT STD_LOGIC;
                    signal AUD_R_from_the_spu : OUT STD_LOGIC;
                    signal DAC_BCLK_from_the_spu : OUT STD_LOGIC;
                    signal DAC_DATA_from_the_spu : OUT STD_LOGIC;
                    signal DAC_LRCK_from_the_spu : OUT STD_LOGIC;
                    signal SPDIF_from_the_spu : OUT STD_LOGIC;
                    signal clk_128fs_to_the_spu : IN STD_LOGIC;

                 -- the_sysuart
                    signal rxd_to_the_sysuart : IN STD_LOGIC;
                    signal txd_from_the_sysuart : OUT STD_LOGIC;

                 -- the_vga
                    signal video_bout_from_the_vga : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal video_clk_to_the_vga : IN STD_LOGIC;
                    signal video_enable_from_the_vga : OUT STD_LOGIC;
                    signal video_gout_from_the_vga : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal video_hsync_n_from_the_vga : OUT STD_LOGIC;
                    signal video_rout_from_the_vga : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal video_vsync_n_from_the_vga : OUT STD_LOGIC
                 );
end component nios2_fpu;

component sdram_test_component is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal zs_addr : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal zs_ba : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_cas_n : IN STD_LOGIC;
                    signal zs_cke : IN STD_LOGIC;
                    signal zs_cs_n : IN STD_LOGIC;
                    signal zs_dqm : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_ras_n : IN STD_LOGIC;
                    signal zs_we_n : IN STD_LOGIC;

                 -- outputs:
                    signal zs_dq : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sdram_test_component;

                signal AUD_L_from_the_spu :  STD_LOGIC;
                signal AUD_R_from_the_spu :  STD_LOGIC;
                signal DAC_BCLK_from_the_spu :  STD_LOGIC;
                signal DAC_DATA_from_the_spu :  STD_LOGIC;
                signal DAC_LRCK_from_the_spu :  STD_LOGIC;
                signal MMC_CD_to_the_mmcdma :  STD_LOGIC;
                signal MMC_SCK_from_the_mmcdma :  STD_LOGIC;
                signal MMC_SDI_to_the_mmcdma :  STD_LOGIC;
                signal MMC_SDO_from_the_mmcdma :  STD_LOGIC;
                signal MMC_WP_to_the_mmcdma :  STD_LOGIC;
                signal MMC_nCS_from_the_mmcdma :  STD_LOGIC;
                signal SPDIF_from_the_spu :  STD_LOGIC;
                signal bidir_port_to_and_from_the_gpio0 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clk :  STD_LOGIC;
                signal clk_128fs_to_the_spu :  STD_LOGIC;
                signal core_clk :  STD_LOGIC;
                signal in_port_to_the_dipsw :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal in_port_to_the_psw :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_a :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fast_fpu_custom_instruction_master_multi_b :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fast_fpu_custom_instruction_master_multi_c :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal nios2_fast_fpu_custom_instruction_master_multi_clk :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_estatus :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_ipending :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fast_fpu_custom_instruction_master_multi_readra :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_readrb :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_reset :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_status :  STD_LOGIC;
                signal nios2_fast_fpu_custom_instruction_master_multi_writerc :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_0_downstream_nativeaddress :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_0_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_1_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_1_downstream_nativeaddress :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_1_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_2_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_2_downstream_nativeaddress :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_3_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_3_downstream_nativeaddress :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal nios2_fpu_burst_3_upstream_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal nios2_fpu_burst_4_downstream_nativeaddress :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_4_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_5_downstream_nativeaddress :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal nios2_fpu_burst_6_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_6_downstream_nativeaddress :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_7_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_burst_7_downstream_nativeaddress :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal nios2_fpu_burst_7_upstream_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal nios2_fpu_burst_8_downstream_debugaccess :  STD_LOGIC;
                signal nios2_fpu_clock_0_in_endofpacket_from_sa :  STD_LOGIC;
                signal out_port_from_the_led :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal peri_clk :  STD_LOGIC;
                signal peripheral_bridge_m1_debugaccess :  STD_LOGIC;
                signal peripheral_bridge_m1_endofpacket :  STD_LOGIC;
                signal reset_n :  STD_LOGIC;
                signal rxd_to_the_sysuart :  STD_LOGIC;
                signal sysid_control_slave_clock :  STD_LOGIC;
                signal sysuart_s1_dataavailable_from_sa :  STD_LOGIC;
                signal sysuart_s1_readyfordata_from_sa :  STD_LOGIC;
                signal txd_from_the_sysuart :  STD_LOGIC;
                signal video_bout_from_the_vga :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal video_clk_to_the_vga :  STD_LOGIC;
                signal video_enable_from_the_vga :  STD_LOGIC;
                signal video_gout_from_the_vga :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal video_hsync_n_from_the_vga :  STD_LOGIC;
                signal video_rout_from_the_vga :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal video_vsync_n_from_the_vga :  STD_LOGIC;
                signal zs_addr_from_the_sdram :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal zs_ba_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal zs_cas_n_from_the_sdram :  STD_LOGIC;
                signal zs_cke_from_the_sdram :  STD_LOGIC;
                signal zs_cs_n_from_the_sdram :  STD_LOGIC;
                signal zs_dq_to_and_from_the_sdram :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal zs_dqm_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal zs_ras_n_from_the_sdram :  STD_LOGIC;
                signal zs_we_n_from_the_sdram :  STD_LOGIC;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your component and signal declaration here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


begin

  --Set us up the Dut
  DUT : nios2_fpu
    port map(
      AUD_L_from_the_spu => AUD_L_from_the_spu,
      AUD_R_from_the_spu => AUD_R_from_the_spu,
      DAC_BCLK_from_the_spu => DAC_BCLK_from_the_spu,
      DAC_DATA_from_the_spu => DAC_DATA_from_the_spu,
      DAC_LRCK_from_the_spu => DAC_LRCK_from_the_spu,
      MMC_SCK_from_the_mmcdma => MMC_SCK_from_the_mmcdma,
      MMC_SDO_from_the_mmcdma => MMC_SDO_from_the_mmcdma,
      MMC_nCS_from_the_mmcdma => MMC_nCS_from_the_mmcdma,
      SPDIF_from_the_spu => SPDIF_from_the_spu,
      bidir_port_to_and_from_the_gpio0 => bidir_port_to_and_from_the_gpio0,
      out_port_from_the_led => out_port_from_the_led,
      txd_from_the_sysuart => txd_from_the_sysuart,
      video_bout_from_the_vga => video_bout_from_the_vga,
      video_enable_from_the_vga => video_enable_from_the_vga,
      video_gout_from_the_vga => video_gout_from_the_vga,
      video_hsync_n_from_the_vga => video_hsync_n_from_the_vga,
      video_rout_from_the_vga => video_rout_from_the_vga,
      video_vsync_n_from_the_vga => video_vsync_n_from_the_vga,
      zs_addr_from_the_sdram => zs_addr_from_the_sdram,
      zs_ba_from_the_sdram => zs_ba_from_the_sdram,
      zs_cas_n_from_the_sdram => zs_cas_n_from_the_sdram,
      zs_cke_from_the_sdram => zs_cke_from_the_sdram,
      zs_cs_n_from_the_sdram => zs_cs_n_from_the_sdram,
      zs_dq_to_and_from_the_sdram => zs_dq_to_and_from_the_sdram,
      zs_dqm_from_the_sdram => zs_dqm_from_the_sdram,
      zs_ras_n_from_the_sdram => zs_ras_n_from_the_sdram,
      zs_we_n_from_the_sdram => zs_we_n_from_the_sdram,
      MMC_CD_to_the_mmcdma => MMC_CD_to_the_mmcdma,
      MMC_SDI_to_the_mmcdma => MMC_SDI_to_the_mmcdma,
      MMC_WP_to_the_mmcdma => MMC_WP_to_the_mmcdma,
      clk_128fs_to_the_spu => clk_128fs_to_the_spu,
      core_clk => core_clk,
      in_port_to_the_dipsw => in_port_to_the_dipsw,
      in_port_to_the_psw => in_port_to_the_psw,
      peri_clk => peri_clk,
      reset_n => reset_n,
      rxd_to_the_sysuart => rxd_to_the_sysuart,
      video_clk_to_the_vga => video_clk_to_the_vga
    );


  --the_sdram_test_component, which is an e_instance
  the_sdram_test_component : sdram_test_component
    port map(
      zs_dq => zs_dq_to_and_from_the_sdram,
      clk => core_clk,
      zs_addr => zs_addr_from_the_sdram,
      zs_ba => zs_ba_from_the_sdram,
      zs_cas_n => zs_cas_n_from_the_sdram,
      zs_cke => zs_cke_from_the_sdram,
      zs_cs_n => zs_cs_n_from_the_sdram,
      zs_dqm => zs_dqm_from_the_sdram,
      zs_ras_n => zs_ras_n_from_the_sdram,
      zs_we_n => zs_we_n_from_the_sdram
    );


  process
  begin
    core_clk <= '0';
    loop
       wait for 4 ns;
       core_clk <= not core_clk;
    end loop;
  end process;
  process
  begin
    peri_clk <= '0';
    loop
       if (peri_clk = '1') then
          wait for 12 ns;
          peri_clk <= not peri_clk;
       else
          wait for 13 ns;
          peri_clk <= not peri_clk;
       end if;
    end loop;
  end process;
  PROCESS
    BEGIN
       reset_n <= '0';
       wait for 80 ns;
       reset_n <= '1'; 
    WAIT;
  END PROCESS;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add additional architecture here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


end europa;



--synthesis translate_on
